`timescale 1ns/1ns
module CSR_PE_tb();
parameter col_length = 8;
parameter word_length = 8;
parameter double_word_length = 16;
parameter kernel_size = 5;
parameter image_size = 28;

reg clk;
reg rst;
reg signed [word_length-1:0] data_in;
reg in_valid;
//reg [6272-1 :0] pe_input_feature_value='hf0_dd_39_f3_f7_06_02_f7_02_f6_fc_15_f9_ff_15_08_fe_fb_f0_01_e5_09_00_f9_1d_fa_f6_ec_fd_f2_fb_f2_eb_f3_fa_f3_12_fc_f8_0b_03_fe_f1_f6_07_f7_eb_0a_17_f5_05_01_18_1f_f1_09_07_04_f3_0c_fa_f6_01_0d_07_e5_06_f8_0e_0b_f9_03_fc_e1_0b_f2_15_fa_0d_ee_08_f9_ed_ff_f8_fc_fa_f8_e8_07_f2_0f_00_da_08_fb_03_06_f2_f0_07_03_06_fb_e9_f5_13_06_fa_0d_05_0a_f1_0d_f6_03_fa_03_17_1c_06_e4_13_03_11_0c_f4_15_fb_0d_fd_07_02_0b_f5_0e_ea_e0_ee_04_f2_fb_01_01_e7_01_ea_07_0e_fc_08_1f_1a_04_fa_ef_02_00_d8_fa_eb_ee_0d_f1_f4_ff_01_fd_18_eb_f2_08_12_04_0b_fb_f7_0a_00_0b_05_f7_f2_0a_1a_e6_15_0e_29_12_f8_08_dd_f9_0f_10_05_df_02_07_f1_fe_01_0c_dc_fb_fb_fb_16_15_e8_f8_02_fe_0e_10_0d_fb_fa_02_fd_e5_03_09_f5_f9_fd_e5_05_0a_03_04_0c_0a_1d_0f_0e_1b_fb_26_f2_ec_08_08_f8_03_08_1b_fc_19_f7_f4_13_00_fc_13_00_1e_12_fc_11_15_11_00_f7_dd_f6_05_0d_f3_1a_13_fd_18_0e_f1_14_09_dd_0a_ed_e6_f1_06_ed_fc_fb_fe_10_07_f0_17_15_03_07_f5_0a_13_06_13_fa_1c_07_05_03_ee_eb_f1_dc_09_f6_fc_fb_04_d9_f9_08_01_08_18_15_25_e6_fe_f9_03_f1_fc_f3_fb_0e_00_f2_f0_0a_f7_06_0b_f8_26_f5_0c_e6_09_f7_fe_fa_04_fa_0b_dc_f8_12_e4_f3_f5_02_0a_f9_20_fd_04_12_fa_fb_03_15_e2_ef_f4_01_19_0c_fd_fc_fc_03_0f_18_f2_05_e9_f2_22_04_ef_f5_03_fd_10_f4_e2_0b_07_02_ec_f8_01_0e_fe_fc_03_ef_eb_f1_f9_04_06_09_15_fc_01_03_f9_0d_ec_f2_2a_e9_01_0b_12_e9_ff_e9_0d_f3_0f_e4_02_08_0d_e9_e3_fc_05_f3_f6_fd_ee_fc_e4_f5_f3_ef_e1_06_f5_0b_00_16_e1_f2_f1_06_03_ff_fa_07_f3_09_f7_0a_0a_0c_ff_1f_f4_0f_ef_fb_15_02_e6_fd_f9_08_f1_ff_f1_eb_11_f4_ea_fd_f3_f0_05_0a_e9_05_0a_f7_e8_f7_f2_11_f4_03_f5_13_e9_fb_fc_04_fb_0a_01_f9_04_00_03_f7_fb_0b_2c_13_0a_10_ec_08_eb_17_fa_1e_05_18_f4_02_01_0a_03_ff_02_f6_f9_f6_00_07_01_01_f2_0d_19_fc_05_ef_f3_0c_e7_0d_e1_07_09_26_ff_f8_0a_cf_f1_e9_08_04_ff_fe_e4_dc_fa_05_fc_23_09_ff_03_09_04_18_1a_f4_02_d7_2a_ed_09_07_14_f0_ff_0f_09_0f_f8_08_f1_21_02_27_fc_f8_fb_ef_11_ee_f9_17_13_01_2c_04_f6_1c_e8_f7_f8_fa_08_13_f6_11_24_fb_00_f4_09_0d_ff_ff_2c_f2_0f_2b_e0_fa_0c_04_25_fa_0a_0c_0c_15_f9_07_f6_fa_f7_07_20_f8_17_10_07_0a_07_1a_04_0b_f6_ff_1a_ef_e6_03_02_06_1f_fb_0c_06_f9_ff_04_1c_ec_f8_09_fc_20_e8_0e_f6_ed_f6_1c_00_e9_f6_07_15_f1_06_12_f9_e7_ef_08_ed_fb_16_fd_13_0d_fa_df_f0_09_e6_fd_f5_09_03_fa_17_fa_2f_16_ff_09_10_04_09_fe_fd_0d_f6_f2_e3_e2_f1_12_1b_ed_fb_18_fe_fd_01_1b_01_01_f3_1d_ff_07_0f_fe_05_ef_ef_38_fc_fb_ee_fc_f0_0e_02_37_0c_f4_1e_e1_04_f4_f4_0a_22_06_01_f0_00_00_1d_0d_fd_1f_f4_06_02_fe_07_ec_12_f7;
reg [6272-1:0] pe_input_feature_value ='hf9_21_00_e9_1c_00_ef_f9_00_00_00_00_05_00_00_14_e4_00_00_00_00_f1_00_00_00_f7_08_00_14_00_00_00_ee_00_00_1b_00_00_00_00_00_e3_df_f4_09_fb_00_00_0d_00_0e_dc_00_00_00_00_00_ea_06_fb_01_00_00_09_13_00_e4_00_00_f1_0b_f4_00_00_00_00_00_fd_00_f3_13_00_01_25_00_05_00_00_fc_00_00_ec_00_fe_00_00_00_00_00_00_00_00_03_f1_00_08_05_00_22_00_00_14_00_04_fd_ff_13_00_00_e2_00_0a_00_fe_00_fc_fa_00_10_00_00_fe_eb_00_00_00_00_f4_00_14_00_f3_1e_07_00_00_00_d7_00_00_10_00_fc_00_ff_00_00_08_00_00_e9_fa_00_00_f0_00_00_04_f4_00_00_00_00_0b_00_10_e9_e8_00_00_f3_00_00_00_08_00_00_e6_00_11_00_00_fa_f6_00_00_00_00_00_0f_f2_00_00_00_fd_fc_00_f1_00_d4_00_0e_00_00_00_00_00_00_00_07_00_0b_01_00_00_00_00_df_00_00_06_00_00_00_00_00_00_01_00_1e_f6_fc_f8_00_00_ef_00_00_00_1b_00_f4_ed_00_00_00_00_00_00_00_00_ff_00_00_00_f5_00_00_00_eb_00_00_00_ef_f5_eb_00_00_00_00_00_0e_00_00_05_11_f4_fb_00_10_00_10_00_f2_00_df_15_00_0d_00_00_f6_f8_08_00_00_00_00_00_00_00_00_00_ec_00_00_13_00_d5_00_00_05_00_00_00_11_00_00_00_00_ef_00_19_00_00_f5_00_00_08_ff_f2_e7_00_00_00_e8_00_fa_00_00_00_e4_08_f2_16_00_00_0e_00_00_00_00_00_00_f9_ec_00_e2_00_00_00_00_00_fb_00_00_1b_02_f1_00_0a_00_1c_fd_00_f9_04_00_e3_0d_00_0c_00_1a_03_df_00_00_00_00_fe_fa_13_00_10_00_00_00_00_f8_00_00_00_00_00_09_00_00_00_00_0c_00_00_00_f8_00_00_fe_00_f3_00_fa_04_0c_00_00_00_00_10_15_f3_00_f4_10_0b_00_1e_ef_00_00_00_f3_00_00_00_00_00_04_00_00_f2_0f_2f_00_00_00_fa_00_00_00_00_10_00_0a_0c_00_ff_00_00_20_ee_00_00_f7_00_00_00_fb_23_08_00_00_00_00_fc_f9_02_00_00_12_00_00_06_00_fc_f8_00_00_00_00_00_f6_f5_00_00_00_ed_01_01_00_00_00_00_f3_00_00_00_06_00_1c_12_00_ee_01_00_00_00_0f_00_00_03_f2_f8_00_00_00_00_00_00_00_fd_e7_00_fd_00_00_00_fa_0a_16_00_dd_00_f1_1e_ef_00_00_00_00_00_00_f5_00_00_00_00_00_00_0f_ef_00_00_00_00_15_1b_00_00_e8_00_00_00_08_00_00_02_00_00_00_00_00_0e_0d_fc_01_02_ff_00_0f_00_00_07_00_00_1f_00_00_00_00_00_00_0f_00_00_0e_e9_00_f3_00_00_00_00_00_00_00_1b_02_00_e1_00_00_00_04_00_00_00_00_00_00_00_06_00_f6_ec_00_0f_07_00_00_f9_01_00_f8_0c_00_00_00_00_00_f8_00_00_00_12_00_00_32_fb_00_00_00_ea_00_00_00_ff_00_e5_00_00_00_00_00_f9_00_00_10_00_00_ec_e4_00_f9_09_00_00_0f_0b_0d_00_12_00_00_fe_ff_00_00_00_14_00_ef_e7_00_00_00_f8_0a_00_00_fe_00_f6_00_00_00_2a_00_00_19_1b_00_fa_00_00_00_f2_00_00_00_00_ed_00_00_f6_f4_00_00_00_00_00_ff_00_00_04_1a_16_03_00_cf_04_00_00_ec_00_02_f6_00_e2_f0_02_00_00_0c;
reg [6272-1 :0] pe_input_feature_rows='h1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1B_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_1A_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_19_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_18_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_17_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_16_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_15_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_14_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_13_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_12_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_11_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0F_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0E_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0D_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0C_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0B_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_0A_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_09_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_08_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_07_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_06_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_05_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_04_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_03_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_02_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;
reg [6272-1 :0] pe_input_feature_cols='h1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00_1B_1A_19_18_17_16_15_14_13_12_11_10_0F_0E_0D_0C_0B_0A_09_08_07_06_05_04_03_02_01_00;
reg [224-1:0] pe_input_weight_value ='hfc_06_02_14_fc_f0_07_12_0c_23_fa_ee_f8_11_12_11_00_0a_d8_15_ff_f6_f1_fd_13;
reg [224-1 :0] pe_input_weight_rows='h04_04_04_04_04_03_03_03_03_03_02_02_02_02_02_01_01_01_01_01_00_00_00_00_00;
reg [224-1 :0] pe_input_weight_cols='h04_03_02_01_00_04_03_02_01_00_04_03_02_01_00_04_03_02_01_00_04_03_02_01_00;

reg [double_word_length-1:0] weight_valid_num='d27;

// CSR wire
wire CSR_valid;
wire [image_size*image_size*word_length-1 :0] CSR_data_out;
wire [image_size*image_size*col_length-1:0] CSR_data_out_cols;
wire [image_size*image_size*col_length-1:0] CSR_data_out_rows;
wire [double_word_length-1:0] valid_num_out;

// PE Wire
reg [double_word_length-1:0] in_channel;
wire [double_word_length-1:0] out_channel;
wire PE_out_valid;
wire [double_word_length-1:0] PE_valid_num;
assign PE_valid_num = 'd784;
wire signed [word_length*2*16 -1:0] PE_data_out;
wire signed [col_length*16 -1:0] PE_data_out_cols;
wire signed [col_length*16 -1:0] PE_data_out_rows;
wire signed [word_length*2-1:0] PE_answer_1_1,PE_answer_1_2,PE_answer_1_3,PE_answer_1_4,PE_answer_2_1,PE_answer_2_2,PE_answer_2_3,PE_answer_2_4;
wire signed [word_length*2-1:0] PE_answer_3_1,PE_answer_3_2,PE_answer_3_3,PE_answer_3_4,PE_answer_4_1,PE_answer_4_2,PE_answer_4_3,PE_answer_4_4; 
wire signed [col_length-1:0] PE_col_answer_1_1,PE_col_answer_1_2,PE_col_answer_1_3,PE_col_answer_1_4,PE_col_answer_2_1,PE_col_answer_2_2,PE_col_answer_2_3,PE_col_answer_2_4,PE_col_answer_3_1,PE_col_answer_3_2,PE_col_answer_3_3,PE_col_answer_3_4,PE_col_answer_4_1,PE_col_answer_4_2,PE_col_answer_4_3,PE_col_answer_4_4; 
wire signed [col_length-1:0] PE_row_answer_1_1,PE_row_answer_1_2,PE_row_answer_1_3,PE_row_answer_1_4,PE_row_answer_2_1,PE_row_answer_2_2,PE_row_answer_2_3,PE_row_answer_2_4,PE_row_answer_3_1,PE_row_answer_3_2,PE_row_answer_3_3,PE_row_answer_3_4,PE_row_answer_4_1,PE_row_answer_4_2,PE_row_answer_4_3,PE_row_answer_4_4; 
assign {PE_col_answer_4_4,PE_col_answer_4_3,PE_col_answer_4_2,PE_col_answer_4_1, PE_col_answer_3_4,PE_col_answer_3_3,PE_col_answer_3_2,PE_col_answer_3_1, PE_col_answer_2_4,PE_col_answer_2_3,PE_col_answer_2_2,PE_col_answer_2_1, PE_col_answer_1_4,PE_col_answer_1_3,PE_col_answer_1_2,PE_col_answer_1_1}= PE_data_out_cols;
assign {PE_row_answer_4_4,PE_row_answer_4_3,PE_row_answer_4_2,PE_row_answer_4_1, PE_row_answer_3_4,PE_row_answer_3_3,PE_row_answer_3_2,PE_row_answer_3_1, PE_row_answer_2_4,PE_row_answer_2_3,PE_row_answer_2_2,PE_row_answer_2_1, PE_row_answer_1_4,PE_row_answer_1_3,PE_row_answer_1_2,PE_row_answer_1_1}= PE_data_out_rows;
assign {{PE_answer_1_4},{PE_answer_1_3},{PE_answer_1_2},{PE_answer_1_1}} = PE_data_out[word_length*2*4 -1 -:word_length*2*4];
assign {{PE_answer_2_4},{PE_answer_2_3},{PE_answer_2_2},{PE_answer_2_1}} = PE_data_out[word_length*2*8 -1 -:word_length*2*4];
assign {{PE_answer_3_4},{PE_answer_3_3},{PE_answer_3_2},{PE_answer_3_1}} = PE_data_out[word_length*2*12 -1 -:word_length*2*4];
assign {{PE_answer_4_4},{PE_answer_4_3},{PE_answer_4_2},{PE_answer_4_1}} = PE_data_out[word_length*2*16 -1 -:word_length*2*4];
reg [32*32*word_length*2-1:0] PE_result;
wire signed  [word_length*2-1:0] PE_pixels_0_0, PE_pixels_0_1, PE_pixels_0_2, PE_pixels_0_3, PE_pixels_0_4, PE_pixels_0_5, PE_pixels_0_6, PE_pixels_0_7, PE_pixels_0_8, PE_pixels_0_9, PE_pixels_0_10, PE_pixels_0_11, PE_pixels_0_12, PE_pixels_0_13, PE_pixels_0_14, PE_pixels_0_15, PE_pixels_0_16, PE_pixels_0_17, PE_pixels_0_18, PE_pixels_0_19, PE_pixels_0_20, PE_pixels_0_21, PE_pixels_0_22, PE_pixels_0_23, PE_pixels_0_24, PE_pixels_0_25, PE_pixels_0_26, PE_pixels_0_27, PE_pixels_0_28, PE_pixels_0_29, PE_pixels_0_30, PE_pixels_0_31, PE_pixels_1_0, PE_pixels_1_1, PE_pixels_1_2, PE_pixels_1_3, PE_pixels_1_4, PE_pixels_1_5, PE_pixels_1_6, PE_pixels_1_7, PE_pixels_1_8, PE_pixels_1_9, PE_pixels_1_10, PE_pixels_1_11, PE_pixels_1_12, PE_pixels_1_13, PE_pixels_1_14, PE_pixels_1_15, PE_pixels_1_16, PE_pixels_1_17, PE_pixels_1_18, PE_pixels_1_19, PE_pixels_1_20, PE_pixels_1_21, PE_pixels_1_22, PE_pixels_1_23, PE_pixels_1_24, PE_pixels_1_25, PE_pixels_1_26, PE_pixels_1_27, PE_pixels_1_28, PE_pixels_1_29, PE_pixels_1_30, PE_pixels_1_31, PE_pixels_2_0, PE_pixels_2_1, PE_pixels_2_2, PE_pixels_2_3, PE_pixels_2_4, PE_pixels_2_5, PE_pixels_2_6, PE_pixels_2_7, PE_pixels_2_8, PE_pixels_2_9, PE_pixels_2_10, PE_pixels_2_11, PE_pixels_2_12, PE_pixels_2_13, PE_pixels_2_14, PE_pixels_2_15, PE_pixels_2_16, PE_pixels_2_17, PE_pixels_2_18, PE_pixels_2_19, PE_pixels_2_20, PE_pixels_2_21, PE_pixels_2_22, PE_pixels_2_23, PE_pixels_2_24, PE_pixels_2_25, PE_pixels_2_26, PE_pixels_2_27, PE_pixels_2_28, PE_pixels_2_29, PE_pixels_2_30, PE_pixels_2_31, PE_pixels_3_0, PE_pixels_3_1, PE_pixels_3_2, PE_pixels_3_3, PE_pixels_3_4, PE_pixels_3_5, PE_pixels_3_6, PE_pixels_3_7, PE_pixels_3_8, PE_pixels_3_9, PE_pixels_3_10, PE_pixels_3_11, PE_pixels_3_12, PE_pixels_3_13, PE_pixels_3_14, PE_pixels_3_15, PE_pixels_3_16, PE_pixels_3_17, PE_pixels_3_18, PE_pixels_3_19, PE_pixels_3_20, PE_pixels_3_21, PE_pixels_3_22, PE_pixels_3_23, PE_pixels_3_24, PE_pixels_3_25, PE_pixels_3_26, PE_pixels_3_27, PE_pixels_3_28, PE_pixels_3_29, PE_pixels_3_30, PE_pixels_3_31, PE_pixels_4_0, PE_pixels_4_1, PE_pixels_4_2, PE_pixels_4_3, PE_pixels_4_4, PE_pixels_4_5, PE_pixels_4_6, PE_pixels_4_7, PE_pixels_4_8, PE_pixels_4_9, PE_pixels_4_10, PE_pixels_4_11, PE_pixels_4_12, PE_pixels_4_13, PE_pixels_4_14, PE_pixels_4_15, PE_pixels_4_16, PE_pixels_4_17, PE_pixels_4_18, PE_pixels_4_19, PE_pixels_4_20, PE_pixels_4_21, PE_pixels_4_22, PE_pixels_4_23, PE_pixels_4_24, PE_pixels_4_25, PE_pixels_4_26, PE_pixels_4_27, PE_pixels_4_28, PE_pixels_4_29, PE_pixels_4_30, PE_pixels_4_31, PE_pixels_5_0, PE_pixels_5_1, PE_pixels_5_2, PE_pixels_5_3, PE_pixels_5_4, PE_pixels_5_5, PE_pixels_5_6, PE_pixels_5_7, PE_pixels_5_8, PE_pixels_5_9, PE_pixels_5_10, PE_pixels_5_11, PE_pixels_5_12, PE_pixels_5_13, PE_pixels_5_14, PE_pixels_5_15, PE_pixels_5_16, PE_pixels_5_17, PE_pixels_5_18, PE_pixels_5_19, PE_pixels_5_20, PE_pixels_5_21, PE_pixels_5_22, PE_pixels_5_23, PE_pixels_5_24, PE_pixels_5_25, PE_pixels_5_26, PE_pixels_5_27, PE_pixels_5_28, PE_pixels_5_29, PE_pixels_5_30, PE_pixels_5_31, PE_pixels_6_0, PE_pixels_6_1, PE_pixels_6_2, PE_pixels_6_3, PE_pixels_6_4, PE_pixels_6_5, PE_pixels_6_6, PE_pixels_6_7, PE_pixels_6_8, PE_pixels_6_9, PE_pixels_6_10, PE_pixels_6_11, PE_pixels_6_12, PE_pixels_6_13, PE_pixels_6_14, PE_pixels_6_15, PE_pixels_6_16, PE_pixels_6_17, PE_pixels_6_18, PE_pixels_6_19, PE_pixels_6_20, PE_pixels_6_21, PE_pixels_6_22, PE_pixels_6_23, PE_pixels_6_24, PE_pixels_6_25, PE_pixels_6_26, PE_pixels_6_27, PE_pixels_6_28, PE_pixels_6_29, PE_pixels_6_30, PE_pixels_6_31, PE_pixels_7_0, PE_pixels_7_1, PE_pixels_7_2, PE_pixels_7_3, PE_pixels_7_4, PE_pixels_7_5, PE_pixels_7_6, PE_pixels_7_7, PE_pixels_7_8, PE_pixels_7_9, PE_pixels_7_10, PE_pixels_7_11, PE_pixels_7_12, PE_pixels_7_13, PE_pixels_7_14, PE_pixels_7_15, PE_pixels_7_16, PE_pixels_7_17, PE_pixels_7_18, PE_pixels_7_19, PE_pixels_7_20, PE_pixels_7_21, PE_pixels_7_22, PE_pixels_7_23, PE_pixels_7_24, PE_pixels_7_25, PE_pixels_7_26, PE_pixels_7_27, PE_pixels_7_28, PE_pixels_7_29, PE_pixels_7_30, PE_pixels_7_31, PE_pixels_8_0, PE_pixels_8_1, PE_pixels_8_2, PE_pixels_8_3, PE_pixels_8_4, PE_pixels_8_5, PE_pixels_8_6, PE_pixels_8_7, PE_pixels_8_8, PE_pixels_8_9, PE_pixels_8_10, PE_pixels_8_11, PE_pixels_8_12, PE_pixels_8_13, PE_pixels_8_14, PE_pixels_8_15, PE_pixels_8_16, PE_pixels_8_17, PE_pixels_8_18, PE_pixels_8_19, PE_pixels_8_20, PE_pixels_8_21, PE_pixels_8_22, PE_pixels_8_23, PE_pixels_8_24, PE_pixels_8_25, PE_pixels_8_26, PE_pixels_8_27, PE_pixels_8_28, PE_pixels_8_29, PE_pixels_8_30, PE_pixels_8_31, PE_pixels_9_0, PE_pixels_9_1, PE_pixels_9_2, PE_pixels_9_3, PE_pixels_9_4, PE_pixels_9_5, PE_pixels_9_6, PE_pixels_9_7, PE_pixels_9_8, PE_pixels_9_9, PE_pixels_9_10, PE_pixels_9_11, PE_pixels_9_12, PE_pixels_9_13, PE_pixels_9_14, PE_pixels_9_15, PE_pixels_9_16, PE_pixels_9_17, PE_pixels_9_18, PE_pixels_9_19, PE_pixels_9_20, PE_pixels_9_21, PE_pixels_9_22, PE_pixels_9_23, PE_pixels_9_24, PE_pixels_9_25, PE_pixels_9_26, PE_pixels_9_27, PE_pixels_9_28, PE_pixels_9_29, PE_pixels_9_30, PE_pixels_9_31, PE_pixels_10_0, PE_pixels_10_1, PE_pixels_10_2, PE_pixels_10_3, PE_pixels_10_4, PE_pixels_10_5, PE_pixels_10_6, PE_pixels_10_7, PE_pixels_10_8, PE_pixels_10_9, PE_pixels_10_10, PE_pixels_10_11, PE_pixels_10_12, PE_pixels_10_13, PE_pixels_10_14, PE_pixels_10_15, PE_pixels_10_16, PE_pixels_10_17, PE_pixels_10_18, PE_pixels_10_19, PE_pixels_10_20, PE_pixels_10_21, PE_pixels_10_22, PE_pixels_10_23, PE_pixels_10_24, PE_pixels_10_25, PE_pixels_10_26, PE_pixels_10_27, PE_pixels_10_28, PE_pixels_10_29, PE_pixels_10_30, PE_pixels_10_31, PE_pixels_11_0, PE_pixels_11_1, PE_pixels_11_2, PE_pixels_11_3, PE_pixels_11_4, PE_pixels_11_5, PE_pixels_11_6, PE_pixels_11_7, PE_pixels_11_8, PE_pixels_11_9, PE_pixels_11_10, PE_pixels_11_11, PE_pixels_11_12, PE_pixels_11_13, PE_pixels_11_14, PE_pixels_11_15, PE_pixels_11_16, PE_pixels_11_17, PE_pixels_11_18, PE_pixels_11_19, PE_pixels_11_20, PE_pixels_11_21, PE_pixels_11_22, PE_pixels_11_23, PE_pixels_11_24, PE_pixels_11_25, PE_pixels_11_26, PE_pixels_11_27, PE_pixels_11_28, PE_pixels_11_29, PE_pixels_11_30, PE_pixels_11_31, PE_pixels_12_0, PE_pixels_12_1, PE_pixels_12_2, PE_pixels_12_3, PE_pixels_12_4, PE_pixels_12_5, PE_pixels_12_6, PE_pixels_12_7, PE_pixels_12_8, PE_pixels_12_9, PE_pixels_12_10, PE_pixels_12_11, PE_pixels_12_12, PE_pixels_12_13, PE_pixels_12_14, PE_pixels_12_15, PE_pixels_12_16, PE_pixels_12_17, PE_pixels_12_18, PE_pixels_12_19, PE_pixels_12_20, PE_pixels_12_21, PE_pixels_12_22, PE_pixels_12_23, PE_pixels_12_24, PE_pixels_12_25, PE_pixels_12_26, PE_pixels_12_27, PE_pixels_12_28, PE_pixels_12_29, PE_pixels_12_30, PE_pixels_12_31, PE_pixels_13_0, PE_pixels_13_1, PE_pixels_13_2, PE_pixels_13_3, PE_pixels_13_4, PE_pixels_13_5, PE_pixels_13_6, PE_pixels_13_7, PE_pixels_13_8, PE_pixels_13_9, PE_pixels_13_10, PE_pixels_13_11, PE_pixels_13_12, PE_pixels_13_13, PE_pixels_13_14, PE_pixels_13_15, PE_pixels_13_16, PE_pixels_13_17, PE_pixels_13_18, PE_pixels_13_19, PE_pixels_13_20, PE_pixels_13_21, PE_pixels_13_22, PE_pixels_13_23, PE_pixels_13_24, PE_pixels_13_25, PE_pixels_13_26, PE_pixels_13_27, PE_pixels_13_28, PE_pixels_13_29, PE_pixels_13_30, PE_pixels_13_31, PE_pixels_14_0, PE_pixels_14_1, PE_pixels_14_2, PE_pixels_14_3, PE_pixels_14_4, PE_pixels_14_5, PE_pixels_14_6, PE_pixels_14_7, PE_pixels_14_8, PE_pixels_14_9, PE_pixels_14_10, PE_pixels_14_11, PE_pixels_14_12, PE_pixels_14_13, PE_pixels_14_14, PE_pixels_14_15, PE_pixels_14_16, PE_pixels_14_17, PE_pixels_14_18, PE_pixels_14_19, PE_pixels_14_20, PE_pixels_14_21, PE_pixels_14_22, PE_pixels_14_23, PE_pixels_14_24, PE_pixels_14_25, PE_pixels_14_26, PE_pixels_14_27, PE_pixels_14_28, PE_pixels_14_29, PE_pixels_14_30, PE_pixels_14_31, PE_pixels_15_0, PE_pixels_15_1, PE_pixels_15_2, PE_pixels_15_3, PE_pixels_15_4, PE_pixels_15_5, PE_pixels_15_6, PE_pixels_15_7, PE_pixels_15_8, PE_pixels_15_9, PE_pixels_15_10, PE_pixels_15_11, PE_pixels_15_12, PE_pixels_15_13, PE_pixels_15_14, PE_pixels_15_15, PE_pixels_15_16, PE_pixels_15_17, PE_pixels_15_18, PE_pixels_15_19, PE_pixels_15_20, PE_pixels_15_21, PE_pixels_15_22, PE_pixels_15_23, PE_pixels_15_24, PE_pixels_15_25, PE_pixels_15_26, PE_pixels_15_27, PE_pixels_15_28, PE_pixels_15_29, PE_pixels_15_30, PE_pixels_15_31, PE_pixels_16_0, PE_pixels_16_1, PE_pixels_16_2, PE_pixels_16_3, PE_pixels_16_4, PE_pixels_16_5, PE_pixels_16_6, PE_pixels_16_7, PE_pixels_16_8, PE_pixels_16_9, PE_pixels_16_10, PE_pixels_16_11, PE_pixels_16_12, PE_pixels_16_13, PE_pixels_16_14, PE_pixels_16_15, PE_pixels_16_16, PE_pixels_16_17, PE_pixels_16_18, PE_pixels_16_19, PE_pixels_16_20, PE_pixels_16_21, PE_pixels_16_22, PE_pixels_16_23, PE_pixels_16_24, PE_pixels_16_25, PE_pixels_16_26, PE_pixels_16_27, PE_pixels_16_28, PE_pixels_16_29, PE_pixels_16_30, PE_pixels_16_31, PE_pixels_17_0, PE_pixels_17_1, PE_pixels_17_2, PE_pixels_17_3, PE_pixels_17_4, PE_pixels_17_5, PE_pixels_17_6, PE_pixels_17_7, PE_pixels_17_8, PE_pixels_17_9, PE_pixels_17_10, PE_pixels_17_11, PE_pixels_17_12, PE_pixels_17_13, PE_pixels_17_14, PE_pixels_17_15, PE_pixels_17_16, PE_pixels_17_17, PE_pixels_17_18, PE_pixels_17_19, PE_pixels_17_20, PE_pixels_17_21, PE_pixels_17_22, PE_pixels_17_23, PE_pixels_17_24, PE_pixels_17_25, PE_pixels_17_26, PE_pixels_17_27, PE_pixels_17_28, PE_pixels_17_29, PE_pixels_17_30, PE_pixels_17_31, PE_pixels_18_0, PE_pixels_18_1, PE_pixels_18_2, PE_pixels_18_3, PE_pixels_18_4, PE_pixels_18_5, PE_pixels_18_6, PE_pixels_18_7, PE_pixels_18_8, PE_pixels_18_9, PE_pixels_18_10, PE_pixels_18_11, PE_pixels_18_12, PE_pixels_18_13, PE_pixels_18_14, PE_pixels_18_15, PE_pixels_18_16, PE_pixels_18_17, PE_pixels_18_18, PE_pixels_18_19, PE_pixels_18_20, PE_pixels_18_21, PE_pixels_18_22, PE_pixels_18_23, PE_pixels_18_24, PE_pixels_18_25, PE_pixels_18_26, PE_pixels_18_27, PE_pixels_18_28, PE_pixels_18_29, PE_pixels_18_30, PE_pixels_18_31, PE_pixels_19_0, PE_pixels_19_1, PE_pixels_19_2, PE_pixels_19_3, PE_pixels_19_4, PE_pixels_19_5, PE_pixels_19_6, PE_pixels_19_7, PE_pixels_19_8, PE_pixels_19_9, PE_pixels_19_10, PE_pixels_19_11, PE_pixels_19_12, PE_pixels_19_13, PE_pixels_19_14, PE_pixels_19_15, PE_pixels_19_16, PE_pixels_19_17, PE_pixels_19_18, PE_pixels_19_19, PE_pixels_19_20, PE_pixels_19_21, PE_pixels_19_22, PE_pixels_19_23, PE_pixels_19_24, PE_pixels_19_25, PE_pixels_19_26, PE_pixels_19_27, PE_pixels_19_28, PE_pixels_19_29, PE_pixels_19_30, PE_pixels_19_31, PE_pixels_20_0, PE_pixels_20_1, PE_pixels_20_2, PE_pixels_20_3, PE_pixels_20_4, PE_pixels_20_5, PE_pixels_20_6, PE_pixels_20_7, PE_pixels_20_8, PE_pixels_20_9, PE_pixels_20_10, PE_pixels_20_11, PE_pixels_20_12, PE_pixels_20_13, PE_pixels_20_14, PE_pixels_20_15, PE_pixels_20_16, PE_pixels_20_17, PE_pixels_20_18, PE_pixels_20_19, PE_pixels_20_20, PE_pixels_20_21, PE_pixels_20_22, PE_pixels_20_23, PE_pixels_20_24, PE_pixels_20_25, PE_pixels_20_26, PE_pixels_20_27, PE_pixels_20_28, PE_pixels_20_29, PE_pixels_20_30, PE_pixels_20_31, PE_pixels_21_0, PE_pixels_21_1, PE_pixels_21_2, PE_pixels_21_3, PE_pixels_21_4, PE_pixels_21_5, PE_pixels_21_6, PE_pixels_21_7, PE_pixels_21_8, PE_pixels_21_9, PE_pixels_21_10, PE_pixels_21_11, PE_pixels_21_12, PE_pixels_21_13, PE_pixels_21_14, PE_pixels_21_15, PE_pixels_21_16, PE_pixels_21_17, PE_pixels_21_18, PE_pixels_21_19, PE_pixels_21_20, PE_pixels_21_21, PE_pixels_21_22, PE_pixels_21_23, PE_pixels_21_24, PE_pixels_21_25, PE_pixels_21_26, PE_pixels_21_27, PE_pixels_21_28, PE_pixels_21_29, PE_pixels_21_30, PE_pixels_21_31, PE_pixels_22_0, PE_pixels_22_1, PE_pixels_22_2, PE_pixels_22_3, PE_pixels_22_4, PE_pixels_22_5, PE_pixels_22_6, PE_pixels_22_7, PE_pixels_22_8, PE_pixels_22_9, PE_pixels_22_10, PE_pixels_22_11, PE_pixels_22_12, PE_pixels_22_13, PE_pixels_22_14, PE_pixels_22_15, PE_pixels_22_16, PE_pixels_22_17, PE_pixels_22_18, PE_pixels_22_19, PE_pixels_22_20, PE_pixels_22_21, PE_pixels_22_22, PE_pixels_22_23, PE_pixels_22_24, PE_pixels_22_25, PE_pixels_22_26, PE_pixels_22_27, PE_pixels_22_28, PE_pixels_22_29, PE_pixels_22_30, PE_pixels_22_31, 
PE_pixels_23_0, PE_pixels_23_1, PE_pixels_23_2, PE_pixels_23_3, PE_pixels_23_4, PE_pixels_23_5, PE_pixels_23_6, PE_pixels_23_7, PE_pixels_23_8, PE_pixels_23_9, PE_pixels_23_10, PE_pixels_23_11, PE_pixels_23_12, PE_pixels_23_13, PE_pixels_23_14, PE_pixels_23_15, PE_pixels_23_16, PE_pixels_23_17, PE_pixels_23_18, PE_pixels_23_19, PE_pixels_23_20, PE_pixels_23_21, PE_pixels_23_22, PE_pixels_23_23, PE_pixels_23_24, PE_pixels_23_25, PE_pixels_23_26, PE_pixels_23_27, PE_pixels_23_28, PE_pixels_23_29, PE_pixels_23_30, PE_pixels_23_31, PE_pixels_24_0, PE_pixels_24_1, PE_pixels_24_2, PE_pixels_24_3, PE_pixels_24_4, PE_pixels_24_5, PE_pixels_24_6, PE_pixels_24_7, PE_pixels_24_8, PE_pixels_24_9, PE_pixels_24_10, PE_pixels_24_11, PE_pixels_24_12, PE_pixels_24_13, PE_pixels_24_14, PE_pixels_24_15, PE_pixels_24_16, PE_pixels_24_17, PE_pixels_24_18, PE_pixels_24_19, PE_pixels_24_20, PE_pixels_24_21, PE_pixels_24_22, PE_pixels_24_23, PE_pixels_24_24, PE_pixels_24_25, PE_pixels_24_26, PE_pixels_24_27, PE_pixels_24_28, PE_pixels_24_29, PE_pixels_24_30, PE_pixels_24_31, PE_pixels_25_0, PE_pixels_25_1, PE_pixels_25_2, PE_pixels_25_3, PE_pixels_25_4, PE_pixels_25_5, PE_pixels_25_6, PE_pixels_25_7, PE_pixels_25_8, PE_pixels_25_9, PE_pixels_25_10, PE_pixels_25_11, PE_pixels_25_12, PE_pixels_25_13, PE_pixels_25_14, PE_pixels_25_15, PE_pixels_25_16, PE_pixels_25_17, PE_pixels_25_18, PE_pixels_25_19, PE_pixels_25_20, PE_pixels_25_21, PE_pixels_25_22, PE_pixels_25_23, PE_pixels_25_24, PE_pixels_25_25, PE_pixels_25_26, PE_pixels_25_27, PE_pixels_25_28, PE_pixels_25_29, PE_pixels_25_30, PE_pixels_25_31, PE_pixels_26_0, PE_pixels_26_1, PE_pixels_26_2, PE_pixels_26_3, PE_pixels_26_4, PE_pixels_26_5, PE_pixels_26_6, PE_pixels_26_7, PE_pixels_26_8, PE_pixels_26_9, PE_pixels_26_10, PE_pixels_26_11, PE_pixels_26_12, PE_pixels_26_13, PE_pixels_26_14, PE_pixels_26_15, PE_pixels_26_16, PE_pixels_26_17, PE_pixels_26_18, PE_pixels_26_19, PE_pixels_26_20, PE_pixels_26_21, PE_pixels_26_22, PE_pixels_26_23, PE_pixels_26_24, PE_pixels_26_25, PE_pixels_26_26, PE_pixels_26_27, PE_pixels_26_28, PE_pixels_26_29, PE_pixels_26_30, PE_pixels_26_31, PE_pixels_27_0, PE_pixels_27_1, PE_pixels_27_2, PE_pixels_27_3, PE_pixels_27_4, PE_pixels_27_5, PE_pixels_27_6, PE_pixels_27_7, PE_pixels_27_8, PE_pixels_27_9, PE_pixels_27_10, PE_pixels_27_11, PE_pixels_27_12, PE_pixels_27_13, PE_pixels_27_14, PE_pixels_27_15, PE_pixels_27_16, PE_pixels_27_17, PE_pixels_27_18, PE_pixels_27_19, PE_pixels_27_20, PE_pixels_27_21, PE_pixels_27_22, PE_pixels_27_23, PE_pixels_27_24, PE_pixels_27_25, PE_pixels_27_26, PE_pixels_27_27, PE_pixels_27_28, PE_pixels_27_29, PE_pixels_27_30, PE_pixels_27_31, PE_pixels_28_0, PE_pixels_28_1, PE_pixels_28_2, PE_pixels_28_3, PE_pixels_28_4, PE_pixels_28_5, PE_pixels_28_6, PE_pixels_28_7, PE_pixels_28_8, PE_pixels_28_9, PE_pixels_28_10, PE_pixels_28_11, PE_pixels_28_12, PE_pixels_28_13, PE_pixels_28_14, PE_pixels_28_15, PE_pixels_28_16, PE_pixels_28_17, PE_pixels_28_18, PE_pixels_28_19, PE_pixels_28_20, PE_pixels_28_21, PE_pixels_28_22, PE_pixels_28_23, PE_pixels_28_24, PE_pixels_28_25, PE_pixels_28_26, PE_pixels_28_27, PE_pixels_28_28, PE_pixels_28_29, PE_pixels_28_30, PE_pixels_28_31, PE_pixels_29_0, PE_pixels_29_1, PE_pixels_29_2, PE_pixels_29_3, PE_pixels_29_4, PE_pixels_29_5, PE_pixels_29_6, PE_pixels_29_7, PE_pixels_29_8, PE_pixels_29_9, PE_pixels_29_10, PE_pixels_29_11, PE_pixels_29_12, PE_pixels_29_13, PE_pixels_29_14, PE_pixels_29_15, PE_pixels_29_16, PE_pixels_29_17, PE_pixels_29_18, PE_pixels_29_19, PE_pixels_29_20, PE_pixels_29_21, PE_pixels_29_22, PE_pixels_29_23, PE_pixels_29_24, PE_pixels_29_25, PE_pixels_29_26, PE_pixels_29_27, PE_pixels_29_28, PE_pixels_29_29, PE_pixels_29_30, PE_pixels_29_31, PE_pixels_30_0, PE_pixels_30_1, PE_pixels_30_2, PE_pixels_30_3, PE_pixels_30_4, PE_pixels_30_5, PE_pixels_30_6, PE_pixels_30_7, PE_pixels_30_8, PE_pixels_30_9, PE_pixels_30_10, PE_pixels_30_11, PE_pixels_30_12, PE_pixels_30_13, PE_pixels_30_14, PE_pixels_30_15, PE_pixels_30_16, PE_pixels_30_17, PE_pixels_30_18, PE_pixels_30_19, PE_pixels_30_20, PE_pixels_30_21, PE_pixels_30_22, PE_pixels_30_23, PE_pixels_30_24, PE_pixels_30_25, PE_pixels_30_26, PE_pixels_30_27, PE_pixels_30_28, PE_pixels_30_29, PE_pixels_30_30, PE_pixels_30_31, PE_pixels_31_0, PE_pixels_31_1, PE_pixels_31_2, PE_pixels_31_3, PE_pixels_31_4, PE_pixels_31_5, PE_pixels_31_6, PE_pixels_31_7, PE_pixels_31_8, PE_pixels_31_9, PE_pixels_31_10, PE_pixels_31_11, PE_pixels_31_12, PE_pixels_31_13, PE_pixels_31_14, PE_pixels_31_15, PE_pixels_31_16, PE_pixels_31_17, PE_pixels_31_18, PE_pixels_31_19, PE_pixels_31_20, PE_pixels_31_21, PE_pixels_31_22, PE_pixels_31_23, PE_pixels_31_24, PE_pixels_31_25, PE_pixels_31_26, PE_pixels_31_27, PE_pixels_31_28, PE_pixels_31_29, PE_pixels_31_30, PE_pixels_31_31;
assign PE_pixels_0_0 = {PE_result[1*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_0 = {PE_result[2*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_0 = {PE_result[3*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_0 = {PE_result[4*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_0 = {PE_result[5*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_0 = {PE_result[6*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_0 = {PE_result[7*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_0 = {PE_result[8*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_0 = {PE_result[9*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_0 = {PE_result[10*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_0 = {PE_result[11*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_0 = {PE_result[12*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_0 = {PE_result[13*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_0 = {PE_result[14*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_0 = {PE_result[15*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_0 = {PE_result[16*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_0 = {PE_result[17*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_0 = {PE_result[18*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_0 = {PE_result[19*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_0 = {PE_result[20*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_0 = {PE_result[21*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_0 = {PE_result[22*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_0 = {PE_result[23*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_0 = {PE_result[24*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_0 = {PE_result[25*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_0 = {PE_result[26*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_0 = {PE_result[27*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_0 = {PE_result[28*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_0 = {PE_result[29*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_0 = {PE_result[30*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_0 = {PE_result[31*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_0 = {PE_result[32*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_1 = {PE_result[33*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_1 = {PE_result[34*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_1 = {PE_result[35*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_1 = {PE_result[36*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_1 = {PE_result[37*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_1 = {PE_result[38*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_1 = {PE_result[39*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_1 = {PE_result[40*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_1 = {PE_result[41*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_1 = {PE_result[42*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_1 = {PE_result[43*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_1 = {PE_result[44*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_1 = {PE_result[45*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_1 = {PE_result[46*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_1 = {PE_result[47*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_1 = {PE_result[48*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_1 = {PE_result[49*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_1 = {PE_result[50*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_1 = {PE_result[51*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_1 = {PE_result[52*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_1 = {PE_result[53*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_1 = {PE_result[54*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_1 = {PE_result[55*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_1 = {PE_result[56*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_1 = {PE_result[57*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_1 = {PE_result[58*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_1 = {PE_result[59*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_1 = {PE_result[60*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_1 = {PE_result[61*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_1 = {PE_result[62*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_1 = {PE_result[63*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_1 = {PE_result[64*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_2 = {PE_result[65*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_2 = {PE_result[66*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_2 = {PE_result[67*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_2 = {PE_result[68*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_2 = {PE_result[69*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_2 = {PE_result[70*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_2 = {PE_result[71*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_2 = {PE_result[72*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_2 = {PE_result[73*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_2 = {PE_result[74*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_2 = {PE_result[75*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_2 = {PE_result[76*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_2 = {PE_result[77*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_2 = {PE_result[78*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_2 = {PE_result[79*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_2 = {PE_result[80*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_2 = {PE_result[81*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_2 = {PE_result[82*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_2 = {PE_result[83*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_2 = {PE_result[84*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_2 = {PE_result[85*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_2 = {PE_result[86*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_2 = {PE_result[87*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_2 = {PE_result[88*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_2 = {PE_result[89*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_2 = {PE_result[90*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_2 = {PE_result[91*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_2 = {PE_result[92*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_2 = {PE_result[93*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_2 = {PE_result[94*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_2 = {PE_result[95*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_2 = {PE_result[96*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_3 = {PE_result[97*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_3 = {PE_result[98*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_3 = {PE_result[99*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_3 = {PE_result[100*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_3 = {PE_result[101*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_3 = {PE_result[102*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_3 = {PE_result[103*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_3 = {PE_result[104*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_3 = {PE_result[105*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_3 = {PE_result[106*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_3 = {PE_result[107*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_3 = {PE_result[108*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_3 = {PE_result[109*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_3 = {PE_result[110*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_3 = {PE_result[111*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_3 = {PE_result[112*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_3 = {PE_result[113*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_3 = {PE_result[114*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_3 = {PE_result[115*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_3 = {PE_result[116*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_3 = {PE_result[117*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_3 = {PE_result[118*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_3 = {PE_result[119*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_3 = {PE_result[120*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_3 = {PE_result[121*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_3 = {PE_result[122*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_3 = {PE_result[123*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_3 = {PE_result[124*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_3 = {PE_result[125*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_3 = {PE_result[126*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_3 = {PE_result[127*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_3 = {PE_result[128*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_4 = {PE_result[129*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_4 = {PE_result[130*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_4 = {PE_result[131*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_4 = {PE_result[132*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_4 = {PE_result[133*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_4 = {PE_result[134*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_4 = {PE_result[135*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_4 = {PE_result[136*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_4 = {PE_result[137*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_4 = {PE_result[138*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_4 = {PE_result[139*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_4 = {PE_result[140*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_4 = {PE_result[141*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_4 = {PE_result[142*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_4 = {PE_result[143*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_4 = {PE_result[144*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_4 = {PE_result[145*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_4 = {PE_result[146*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_4 = {PE_result[147*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_4 = {PE_result[148*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_4 = {PE_result[149*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_4 = {PE_result[150*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_4 = {PE_result[151*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_4 = {PE_result[152*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_4 = {PE_result[153*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_4 = {PE_result[154*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_4 = {PE_result[155*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_4 = {PE_result[156*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_4 = {PE_result[157*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_4 = {PE_result[158*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_4 = {PE_result[159*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_4 = {PE_result[160*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_5 = {PE_result[161*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_5 = {PE_result[162*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_5 = {PE_result[163*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_5 = {PE_result[164*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_5 = {PE_result[165*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_5 = {PE_result[166*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_5 = {PE_result[167*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_5 = {PE_result[168*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_5 = {PE_result[169*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_5 = {PE_result[170*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_5 = {PE_result[171*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_5 = {PE_result[172*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_5 = {PE_result[173*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_5 = {PE_result[174*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_5 = {PE_result[175*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_5 = {PE_result[176*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_5 = {PE_result[177*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_5 = {PE_result[178*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_5 = {PE_result[179*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_5 = {PE_result[180*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_5 = {PE_result[181*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_5 = {PE_result[182*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_5 = {PE_result[183*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_5 = {PE_result[184*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_5 = {PE_result[185*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_5 = {PE_result[186*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_5 = {PE_result[187*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_5 = {PE_result[188*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_5 = {PE_result[189*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_5 = {PE_result[190*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_5 = {PE_result[191*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_5 = {PE_result[192*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_6 = {PE_result[193*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_6 = {PE_result[194*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_6 = {PE_result[195*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_6 = {PE_result[196*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_6 = {PE_result[197*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_6 = {PE_result[198*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_6 = {PE_result[199*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_6 = {PE_result[200*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_6 = {PE_result[201*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_6 = {PE_result[202*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_6 = {PE_result[203*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_6 = {PE_result[204*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_6 = {PE_result[205*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_6 = {PE_result[206*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_6 = {PE_result[207*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_6 = {PE_result[208*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_6 = {PE_result[209*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_6 = {PE_result[210*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_6 = {PE_result[211*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_6 = {PE_result[212*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_6 = {PE_result[213*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_6 = {PE_result[214*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_6 = {PE_result[215*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_6 = {PE_result[216*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_6 = {PE_result[217*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_6 = {PE_result[218*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_6 = {PE_result[219*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_6 = {PE_result[220*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_6 = {PE_result[221*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_6 = {PE_result[222*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_6 = {PE_result[223*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_6 = {PE_result[224*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_7 = {PE_result[225*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_7 = {PE_result[226*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_7 = {PE_result[227*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_7 = {PE_result[228*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_7 = {PE_result[229*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_7 = {PE_result[230*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_7 = {PE_result[231*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_7 = {PE_result[232*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_7 = {PE_result[233*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_7 = {PE_result[234*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_7 = {PE_result[235*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_7 = {PE_result[236*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_7 = {PE_result[237*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_7 = {PE_result[238*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_7 = {PE_result[239*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_7 = {PE_result[240*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_7 = {PE_result[241*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_7 = {PE_result[242*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_7 = {PE_result[243*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_7 = {PE_result[244*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_7 = {PE_result[245*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_7 = {PE_result[246*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_7 = {PE_result[247*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_7 = {PE_result[248*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_7 = {PE_result[249*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_7 = {PE_result[250*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_7 = {PE_result[251*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_7 = {PE_result[252*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_7 = {PE_result[253*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_7 = {PE_result[254*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_7 = {PE_result[255*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_7 = {PE_result[256*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_8 = {PE_result[257*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_8 = {PE_result[258*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_8 = {PE_result[259*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_8 = {PE_result[260*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_8 = {PE_result[261*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_8 = {PE_result[262*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_8 = {PE_result[263*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_8 = {PE_result[264*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_8 = {PE_result[265*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_8 = {PE_result[266*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_8 = {PE_result[267*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_8 = {PE_result[268*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_8 = {PE_result[269*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_8 = {PE_result[270*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_8 = {PE_result[271*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_8 = {PE_result[272*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_8 = {PE_result[273*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_8 = {PE_result[274*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_8 = {PE_result[275*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_8 = {PE_result[276*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_8 = {PE_result[277*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_8 = {PE_result[278*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_8 = {PE_result[279*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_8 = {PE_result[280*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_8 = {PE_result[281*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_8 = {PE_result[282*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_8 = {PE_result[283*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_8 = {PE_result[284*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_8 = {PE_result[285*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_8 = {PE_result[286*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_8 = {PE_result[287*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_8 = {PE_result[288*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_9 = {PE_result[289*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_9 = {PE_result[290*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_9 = {PE_result[291*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_9 = {PE_result[292*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_9 = {PE_result[293*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_9 = {PE_result[294*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_9 = {PE_result[295*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_9 = {PE_result[296*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_9 = {PE_result[297*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_9 = {PE_result[298*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_9 = {PE_result[299*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_9 = {PE_result[300*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_9 = {PE_result[301*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_9 = {PE_result[302*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_9 = {PE_result[303*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_9 = {PE_result[304*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_9 = {PE_result[305*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_9 = {PE_result[306*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_9 = {PE_result[307*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_9 = {PE_result[308*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_9 = {PE_result[309*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_9 = {PE_result[310*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_9 = {PE_result[311*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_9 = {PE_result[312*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_9 = {PE_result[313*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_9 = {PE_result[314*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_9 = {PE_result[315*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_9 = {PE_result[316*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_9 = {PE_result[317*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_9 = {PE_result[318*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_9 = {PE_result[319*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_9 = {PE_result[320*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_10 = {PE_result[321*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_10 = {PE_result[322*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_10 = {PE_result[323*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_10 = {PE_result[324*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_10 = {PE_result[325*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_10 = {PE_result[326*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_10 = {PE_result[327*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_10 = {PE_result[328*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_10 = {PE_result[329*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_10 = {PE_result[330*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_10 = {PE_result[331*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_10 = {PE_result[332*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_10 = {PE_result[333*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_10 = {PE_result[334*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_10 = {PE_result[335*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_10 = {PE_result[336*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_10 = {PE_result[337*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_10 = {PE_result[338*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_10 = {PE_result[339*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_10 = {PE_result[340*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_10 = {PE_result[341*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_10 = {PE_result[342*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_10 = {PE_result[343*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_10 = {PE_result[344*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_10 = {PE_result[345*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_10 = {PE_result[346*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_10 = {PE_result[347*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_10 = {PE_result[348*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_10 = {PE_result[349*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_10 = {PE_result[350*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_10 = {PE_result[351*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_10 = {PE_result[352*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_11 = {PE_result[353*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_11 = {PE_result[354*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_11 = {PE_result[355*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_11 = {PE_result[356*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_11 = {PE_result[357*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_11 = {PE_result[358*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_11 = {PE_result[359*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_11 = {PE_result[360*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_11 = {PE_result[361*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_11 = {PE_result[362*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_11 = {PE_result[363*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_11 = {PE_result[364*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_11 = {PE_result[365*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_11 = {PE_result[366*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_11 = {PE_result[367*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_11 = {PE_result[368*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_11 = {PE_result[369*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_11 = {PE_result[370*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_11 = {PE_result[371*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_11 = {PE_result[372*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_11 = {PE_result[373*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_11 = {PE_result[374*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_11 = {PE_result[375*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_11 = {PE_result[376*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_11 = {PE_result[377*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_11 = {PE_result[378*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_11 = {PE_result[379*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_11 = {PE_result[380*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_11 = {PE_result[381*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_11 = {PE_result[382*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_11 = {PE_result[383*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_11 = {PE_result[384*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_12 = {PE_result[385*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_12 = {PE_result[386*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_12 = {PE_result[387*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_12 = {PE_result[388*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_12 = {PE_result[389*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_12 = {PE_result[390*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_12 = {PE_result[391*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_12 = {PE_result[392*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_12 = {PE_result[393*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_12 = {PE_result[394*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_12 = {PE_result[395*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_12 = {PE_result[396*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_12 = {PE_result[397*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_12 = {PE_result[398*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_12 = {PE_result[399*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_12 = {PE_result[400*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_12 = {PE_result[401*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_12 = {PE_result[402*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_12 = {PE_result[403*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_12 = {PE_result[404*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_12 = {PE_result[405*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_12 = {PE_result[406*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_12 = {PE_result[407*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_12 = {PE_result[408*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_12 = {PE_result[409*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_12 = {PE_result[410*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_12 = {PE_result[411*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_12 = {PE_result[412*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_12 = {PE_result[413*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_12 = {PE_result[414*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_12 = {PE_result[415*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_12 = {PE_result[416*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_13 = {PE_result[417*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_13 = {PE_result[418*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_13 = {PE_result[419*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_13 = {PE_result[420*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_13 = {PE_result[421*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_13 = {PE_result[422*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_13 = {PE_result[423*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_13 = {PE_result[424*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_13 = {PE_result[425*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_13 = {PE_result[426*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_13 = {PE_result[427*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_13 = {PE_result[428*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_13 = {PE_result[429*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_13 = {PE_result[430*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_13 = {PE_result[431*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_13 = {PE_result[432*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_13 = {PE_result[433*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_13 = {PE_result[434*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_13 = {PE_result[435*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_13 = {PE_result[436*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_13 = {PE_result[437*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_13 = {PE_result[438*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_13 = {PE_result[439*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_13 = {PE_result[440*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_13 = {PE_result[441*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_13 = {PE_result[442*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_13 = {PE_result[443*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_13 = {PE_result[444*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_13 = {PE_result[445*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_13 = {PE_result[446*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_13 = {PE_result[447*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_13 = {PE_result[448*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_14 = {PE_result[449*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_14 = {PE_result[450*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_14 = {PE_result[451*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_14 = {PE_result[452*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_14 = {PE_result[453*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_14 = {PE_result[454*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_14 = {PE_result[455*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_14 = {PE_result[456*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_14 = {PE_result[457*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_14 = {PE_result[458*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_14 = {PE_result[459*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_14 = {PE_result[460*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_14 = {PE_result[461*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_14 = {PE_result[462*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_14 = {PE_result[463*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_14 = {PE_result[464*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_14 = {PE_result[465*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_14 = {PE_result[466*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_14 = {PE_result[467*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_14 = {PE_result[468*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_14 = {PE_result[469*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_14 = {PE_result[470*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_14 = {PE_result[471*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_14 = {PE_result[472*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_14 = {PE_result[473*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_14 = {PE_result[474*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_14 = {PE_result[475*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_14 = {PE_result[476*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_14 = {PE_result[477*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_14 = {PE_result[478*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_14 = {PE_result[479*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_14 = {PE_result[480*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_15 = {PE_result[481*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_15 = {PE_result[482*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_15 = {PE_result[483*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_15 = {PE_result[484*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_15 = {PE_result[485*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_15 = {PE_result[486*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_15 = {PE_result[487*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_15 = {PE_result[488*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_15 = {PE_result[489*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_15 = {PE_result[490*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_15 = {PE_result[491*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_15 = {PE_result[492*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_15 = {PE_result[493*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_15 = {PE_result[494*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_15 = {PE_result[495*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_15 = {PE_result[496*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_15 = {PE_result[497*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_15 = {PE_result[498*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_15 = {PE_result[499*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_15 = {PE_result[500*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_15 = {PE_result[501*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_15 = {PE_result[502*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_15 = {PE_result[503*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_15 = {PE_result[504*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_15 = {PE_result[505*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_15 = {PE_result[506*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_15 = {PE_result[507*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_15 = {PE_result[508*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_15 = {PE_result[509*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_15 = {PE_result[510*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_15 = {PE_result[511*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_15 = {PE_result[512*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_16 = {PE_result[513*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_16 = {PE_result[514*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_16 = {PE_result[515*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_16 = {PE_result[516*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_16 = {PE_result[517*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_16 = {PE_result[518*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_16 = {PE_result[519*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_16 = {PE_result[520*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_16 = {PE_result[521*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_16 = {PE_result[522*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_16 = {PE_result[523*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_16 = {PE_result[524*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_16 = {PE_result[525*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_16 = {PE_result[526*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_16 = {PE_result[527*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_16 = {PE_result[528*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_16 = {PE_result[529*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_16 = {PE_result[530*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_16 = {PE_result[531*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_16 = {PE_result[532*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_16 = {PE_result[533*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_16 = {PE_result[534*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_16 = {PE_result[535*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_16 = {PE_result[536*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_16 = {PE_result[537*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_16 = {PE_result[538*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_16 = {PE_result[539*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_16 = {PE_result[540*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_16 = {PE_result[541*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_16 = {PE_result[542*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_16 = {PE_result[543*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_16 = {PE_result[544*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_17 = {PE_result[545*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_17 = {PE_result[546*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_17 = {PE_result[547*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_17 = {PE_result[548*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_17 = {PE_result[549*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_17 = {PE_result[550*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_17 = {PE_result[551*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_17 = {PE_result[552*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_17 = {PE_result[553*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_17 = {PE_result[554*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_17 = {PE_result[555*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_17 = {PE_result[556*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_17 = {PE_result[557*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_17 = {PE_result[558*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_17 = {PE_result[559*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_17 = {PE_result[560*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_17 = {PE_result[561*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_17 = {PE_result[562*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_17 = {PE_result[563*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_17 = {PE_result[564*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_17 = {PE_result[565*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_17 = {PE_result[566*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_17 = {PE_result[567*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_17 = {PE_result[568*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_17 = {PE_result[569*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_17 = {PE_result[570*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_17 = {PE_result[571*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_17 = {PE_result[572*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_17 = {PE_result[573*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_17 = {PE_result[574*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_17 = {PE_result[575*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_17 = {PE_result[576*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_18 = {PE_result[577*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_18 = {PE_result[578*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_18 = {PE_result[579*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_18 = {PE_result[580*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_18 = {PE_result[581*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_18 = {PE_result[582*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_18 = {PE_result[583*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_18 = {PE_result[584*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_18 = {PE_result[585*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_18 = {PE_result[586*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_18 = {PE_result[587*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_18 = {PE_result[588*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_18 = {PE_result[589*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_18 = {PE_result[590*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_18 = {PE_result[591*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_18 = {PE_result[592*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_18 = {PE_result[593*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_18 = {PE_result[594*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_18 = {PE_result[595*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_18 = {PE_result[596*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_18 = {PE_result[597*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_18 = {PE_result[598*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_18 = {PE_result[599*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_18 = {PE_result[600*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_18 = {PE_result[601*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_18 = {PE_result[602*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_18 = {PE_result[603*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_18 = {PE_result[604*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_18 = {PE_result[605*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_18 = {PE_result[606*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_18 = {PE_result[607*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_18 = {PE_result[608*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_19 = {PE_result[609*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_19 = {PE_result[610*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_19 = {PE_result[611*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_19 = {PE_result[612*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_19 = {PE_result[613*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_19 = {PE_result[614*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_19 = {PE_result[615*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_19 = {PE_result[616*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_19 = {PE_result[617*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_19 = {PE_result[618*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_19 = {PE_result[619*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_19 = {PE_result[620*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_19 = {PE_result[621*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_19 = {PE_result[622*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_19 = {PE_result[623*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_19 = {PE_result[624*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_19 = {PE_result[625*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_19 = {PE_result[626*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_19 = {PE_result[627*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_19 = {PE_result[628*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_19 = {PE_result[629*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_19 = {PE_result[630*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_19 = {PE_result[631*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_19 = {PE_result[632*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_19 = {PE_result[633*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_19 = {PE_result[634*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_19 = {PE_result[635*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_19 = {PE_result[636*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_19 = {PE_result[637*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_19 = {PE_result[638*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_19 = {PE_result[639*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_19 = {PE_result[640*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_20 = {PE_result[641*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_20 = {PE_result[642*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_20 = {PE_result[643*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_20 = {PE_result[644*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_20 = {PE_result[645*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_20 = {PE_result[646*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_20 = {PE_result[647*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_20 = {PE_result[648*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_20 = {PE_result[649*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_20 = {PE_result[650*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_20 = {PE_result[651*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_20 = {PE_result[652*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_20 = {PE_result[653*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_20 = {PE_result[654*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_20 = {PE_result[655*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_20 = {PE_result[656*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_20 = {PE_result[657*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_20 = {PE_result[658*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_20 = {PE_result[659*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_20 = {PE_result[660*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_20 = {PE_result[661*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_20 = {PE_result[662*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_20 = {PE_result[663*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_20 = {PE_result[664*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_20 = {PE_result[665*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_20 = {PE_result[666*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_20 = {PE_result[667*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_20 = {PE_result[668*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_20 = {PE_result[669*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_20 = {PE_result[670*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_20 = {PE_result[671*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_20 = {PE_result[672*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_21 = {PE_result[673*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_21 = {PE_result[674*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_21 = {PE_result[675*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_21 = {PE_result[676*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_21 = {PE_result[677*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_21 = {PE_result[678*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_21 = {PE_result[679*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_21 = {PE_result[680*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_21 = {PE_result[681*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_21 = {PE_result[682*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_21 = {PE_result[683*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_21 = {PE_result[684*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_21 = {PE_result[685*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_21 = {PE_result[686*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_21 = {PE_result[687*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_21 = {PE_result[688*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_21 = {PE_result[689*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_21 = {PE_result[690*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_21 = {PE_result[691*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_21 = {PE_result[692*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_21 = {PE_result[693*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_21 = {PE_result[694*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_21 = {PE_result[695*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_21 = {PE_result[696*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_21 = {PE_result[697*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_21 = {PE_result[698*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_21 = {PE_result[699*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_21 = {PE_result[700*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_21 = {PE_result[701*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_21 = {PE_result[702*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_21 = {PE_result[703*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_21 = {PE_result[704*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_22 = {PE_result[705*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_22 = {PE_result[706*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_22 = {PE_result[707*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_22 = {PE_result[708*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_22 = {PE_result[709*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_22 = {PE_result[710*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_22 = {PE_result[711*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_22 = {PE_result[712*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_22 = {PE_result[713*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_22 = {PE_result[714*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_22 = {PE_result[715*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_22 = {PE_result[716*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_22 = {PE_result[717*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_22 = {PE_result[718*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_22 = {PE_result[719*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_22 = {PE_result[720*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_22 = {PE_result[721*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_22 = {PE_result[722*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_22 = {PE_result[723*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_22 = {PE_result[724*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_22 = {PE_result[725*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_22 = {PE_result[726*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_22 = {PE_result[727*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_22 = {PE_result[728*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_22 = {PE_result[729*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_22 = {PE_result[730*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_22 = {PE_result[731*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_22 = {PE_result[732*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_22 = {PE_result[733*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_22 = {PE_result[734*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_22 = {PE_result[735*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_22 = {PE_result[736*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_23 = {PE_result[737*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_23 = {PE_result[738*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_23 = {PE_result[739*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_23 = {PE_result[740*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_23 = {PE_result[741*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_23 = {PE_result[742*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_23 = {PE_result[743*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_23 = {PE_result[744*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_23 = {PE_result[745*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_23 = {PE_result[746*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_23 = {PE_result[747*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_23 = {PE_result[748*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_23 = {PE_result[749*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_23 = {PE_result[750*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_23 = {PE_result[751*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_23 = {PE_result[752*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_23 = {PE_result[753*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_23 = {PE_result[754*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_23 = {PE_result[755*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_23 = {PE_result[756*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_23 = {PE_result[757*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_23 = {PE_result[758*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_23 = {PE_result[759*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_23 = {PE_result[760*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_23 = {PE_result[761*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_23 = {PE_result[762*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_23 = {PE_result[763*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_23 = {PE_result[764*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_23 = {PE_result[765*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_23 = {PE_result[766*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_23 = {PE_result[767*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_23 = {PE_result[768*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_24 = {PE_result[769*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_24 = {PE_result[770*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_24 = {PE_result[771*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_24 = {PE_result[772*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_24 = {PE_result[773*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_24 = {PE_result[774*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_24 = {PE_result[775*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_24 = {PE_result[776*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_24 = {PE_result[777*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_24 = {PE_result[778*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_24 = {PE_result[779*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_24 = {PE_result[780*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_24 = {PE_result[781*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_24 = {PE_result[782*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_24 = {PE_result[783*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_24 = {PE_result[784*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_24 = {PE_result[785*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_24 = {PE_result[786*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_24 = {PE_result[787*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_24 = {PE_result[788*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_24 = {PE_result[789*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_24 = {PE_result[790*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_24 = {PE_result[791*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_24 = {PE_result[792*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_24 = {PE_result[793*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_24 = {PE_result[794*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_24 = {PE_result[795*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_24 = {PE_result[796*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_24 = {PE_result[797*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_24 = {PE_result[798*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_24 = {PE_result[799*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_24 = {PE_result[800*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_25 = {PE_result[801*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_25 = {PE_result[802*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_25 = {PE_result[803*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_25 = {PE_result[804*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_25 = {PE_result[805*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_25 = {PE_result[806*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_25 = {PE_result[807*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_25 = {PE_result[808*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_25 = {PE_result[809*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_25 = {PE_result[810*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_25 = {PE_result[811*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_25 = {PE_result[812*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_25 = {PE_result[813*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_25 = {PE_result[814*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_25 = {PE_result[815*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_25 = {PE_result[816*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_25 = {PE_result[817*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_25 = {PE_result[818*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_25 = {PE_result[819*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_25 = {PE_result[820*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_25 = {PE_result[821*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_25 = {PE_result[822*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_25 = {PE_result[823*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_25 = {PE_result[824*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_25 = {PE_result[825*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_25 = {PE_result[826*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_25 = {PE_result[827*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_25 = {PE_result[828*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_25 = {PE_result[829*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_25 = {PE_result[830*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_25 = {PE_result[831*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_25 = {PE_result[832*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_26 = {PE_result[833*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_26 = {PE_result[834*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_26 = {PE_result[835*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_26 = {PE_result[836*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_26 = {PE_result[837*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_26 = {PE_result[838*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_26 = {PE_result[839*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_26 = {PE_result[840*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_26 = {PE_result[841*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_26 = {PE_result[842*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_26 = {PE_result[843*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_26 = {PE_result[844*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_26 = {PE_result[845*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_26 = {PE_result[846*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_26 = {PE_result[847*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_26 = {PE_result[848*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_26 = {PE_result[849*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_26 = {PE_result[850*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_26 = {PE_result[851*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_26 = {PE_result[852*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_26 = {PE_result[853*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_26 = {PE_result[854*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_26 = {PE_result[855*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_26 = {PE_result[856*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_26 = {PE_result[857*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_26 = {PE_result[858*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_26 = {PE_result[859*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_26 = {PE_result[860*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_26 = {PE_result[861*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_26 = {PE_result[862*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_26 = {PE_result[863*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_26 = {PE_result[864*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_27 = {PE_result[865*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_27 = {PE_result[866*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_27 = {PE_result[867*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_27 = {PE_result[868*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_27 = {PE_result[869*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_27 = {PE_result[870*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_27 = {PE_result[871*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_27 = {PE_result[872*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_27 = {PE_result[873*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_27 = {PE_result[874*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_27 = {PE_result[875*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_27 = {PE_result[876*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_27 = {PE_result[877*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_27 = {PE_result[878*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_27 = {PE_result[879*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_27 = {PE_result[880*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_27 = {PE_result[881*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_27 = {PE_result[882*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_27 = {PE_result[883*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_27 = {PE_result[884*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_27 = {PE_result[885*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_27 = {PE_result[886*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_27 = {PE_result[887*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_27 = {PE_result[888*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_27 = {PE_result[889*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_27 = {PE_result[890*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_27 = {PE_result[891*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_27 = {PE_result[892*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_27 = {PE_result[893*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_27 = {PE_result[894*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_27 = {PE_result[895*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_27 = {PE_result[896*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_28 = {PE_result[897*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_28 = {PE_result[898*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_28 = {PE_result[899*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_28 = {PE_result[900*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_28 = {PE_result[901*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_28 = {PE_result[902*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_28 = {PE_result[903*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_28 = {PE_result[904*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_28 = {PE_result[905*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_28 = {PE_result[906*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_28 = {PE_result[907*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_28 = {PE_result[908*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_28 = {PE_result[909*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_28 = {PE_result[910*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_28 = {PE_result[911*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_28 = {PE_result[912*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_28 = {PE_result[913*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_28 = {PE_result[914*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_28 = {PE_result[915*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_28 = {PE_result[916*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_28 = {PE_result[917*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_28 = {PE_result[918*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_28 = {PE_result[919*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_28 = {PE_result[920*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_28 = {PE_result[921*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_28 = {PE_result[922*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_28 = {PE_result[923*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_28 = {PE_result[924*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_28 = {PE_result[925*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_28 = {PE_result[926*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_28 = {PE_result[927*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_28 = {PE_result[928*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_29 = {PE_result[929*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_29 = {PE_result[930*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_29 = {PE_result[931*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_29 = {PE_result[932*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_29 = {PE_result[933*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_29 = {PE_result[934*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_29 = {PE_result[935*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_29 = {PE_result[936*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_29 = {PE_result[937*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_29 = {PE_result[938*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_29 = {PE_result[939*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_29 = {PE_result[940*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_29 = {PE_result[941*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_29 = {PE_result[942*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_29 = {PE_result[943*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_29 = {PE_result[944*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_29 = {PE_result[945*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_29 = {PE_result[946*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_29 = {PE_result[947*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_29 = {PE_result[948*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_29 = {PE_result[949*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_29 = {PE_result[950*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_29 = {PE_result[951*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_29 = {PE_result[952*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_29 = {PE_result[953*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_29 = {PE_result[954*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_29 = {PE_result[955*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_29 = {PE_result[956*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_29 = {PE_result[957*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_29 = {PE_result[958*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_29 = {PE_result[959*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_29 = {PE_result[960*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_30 = {PE_result[961*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_30 = {PE_result[962*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_30 = {PE_result[963*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_30 = {PE_result[964*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_30 = {PE_result[965*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_30 = {PE_result[966*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_30 = {PE_result[967*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_30 = {PE_result[968*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_30 = {PE_result[969*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_30 = {PE_result[970*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_30 = {PE_result[971*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_30 = {PE_result[972*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_30 = {PE_result[973*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_30 = {PE_result[974*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_30 = {PE_result[975*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_30 = {PE_result[976*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_30 = {PE_result[977*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_30 = {PE_result[978*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_30 = {PE_result[979*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_30 = {PE_result[980*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_30 = {PE_result[981*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_30 = {PE_result[982*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_30 = {PE_result[983*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_30 = {PE_result[984*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_30 = {PE_result[985*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_30 = {PE_result[986*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_30 = {PE_result[987*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_30 = {PE_result[988*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_30 = {PE_result[989*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_30 = {PE_result[990*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_30 = {PE_result[991*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_30 = {PE_result[992*word_length*2-1 -: word_length*2]};
assign PE_pixels_0_31 = {PE_result[993*word_length*2-1 -: word_length*2]};
assign PE_pixels_1_31 = {PE_result[994*word_length*2-1 -: word_length*2]};
assign PE_pixels_2_31 = {PE_result[995*word_length*2-1 -: word_length*2]};
assign PE_pixels_3_31 = {PE_result[996*word_length*2-1 -: word_length*2]};
assign PE_pixels_4_31 = {PE_result[997*word_length*2-1 -: word_length*2]};
assign PE_pixels_5_31 = {PE_result[998*word_length*2-1 -: word_length*2]};
assign PE_pixels_6_31 = {PE_result[999*word_length*2-1 -: word_length*2]};
assign PE_pixels_7_31 = {PE_result[1000*word_length*2-1 -: word_length*2]};
assign PE_pixels_8_31 = {PE_result[1001*word_length*2-1 -: word_length*2]};
assign PE_pixels_9_31 = {PE_result[1002*word_length*2-1 -: word_length*2]};
assign PE_pixels_10_31 = {PE_result[1003*word_length*2-1 -: word_length*2]};
assign PE_pixels_11_31 = {PE_result[1004*word_length*2-1 -: word_length*2]};
assign PE_pixels_12_31 = {PE_result[1005*word_length*2-1 -: word_length*2]};
assign PE_pixels_13_31 = {PE_result[1006*word_length*2-1 -: word_length*2]};
assign PE_pixels_14_31 = {PE_result[1007*word_length*2-1 -: word_length*2]};
assign PE_pixels_15_31 = {PE_result[1008*word_length*2-1 -: word_length*2]};
assign PE_pixels_16_31 = {PE_result[1009*word_length*2-1 -: word_length*2]};
assign PE_pixels_17_31 = {PE_result[1010*word_length*2-1 -: word_length*2]};
assign PE_pixels_18_31 = {PE_result[1011*word_length*2-1 -: word_length*2]};
assign PE_pixels_19_31 = {PE_result[1012*word_length*2-1 -: word_length*2]};
assign PE_pixels_20_31 = {PE_result[1013*word_length*2-1 -: word_length*2]};
assign PE_pixels_21_31 = {PE_result[1014*word_length*2-1 -: word_length*2]};
assign PE_pixels_22_31 = {PE_result[1015*word_length*2-1 -: word_length*2]};
assign PE_pixels_23_31 = {PE_result[1016*word_length*2-1 -: word_length*2]};
assign PE_pixels_24_31 = {PE_result[1017*word_length*2-1 -: word_length*2]};
assign PE_pixels_25_31 = {PE_result[1018*word_length*2-1 -: word_length*2]};
assign PE_pixels_26_31 = {PE_result[1019*word_length*2-1 -: word_length*2]};
assign PE_pixels_27_31 = {PE_result[1020*word_length*2-1 -: word_length*2]};
assign PE_pixels_28_31 = {PE_result[1021*word_length*2-1 -: word_length*2]};
assign PE_pixels_29_31 = {PE_result[1022*word_length*2-1 -: word_length*2]};
assign PE_pixels_30_31 = {PE_result[1023*word_length*2-1 -: word_length*2]};
assign PE_pixels_31_31 = {PE_result[1024*word_length*2-1 -: word_length*2]};

//iter
integer i;
initial begin
    #0      rst = 0;
            clk = 1;
            PE_result = 0;
            data_in = 0;
            in_valid = 0;
            in_channel = 'd1;
    #10     rst = 1;
    #10     rst = 0;
    #100    in_valid = 1;
            for (i=0;i<(image_size*image_size);i=i+1)begin
                data_in[word_length-1:0] = {pe_input_feature_value[(i+1)*word_length-1 -:word_length]};
                #10;
            end
    while(!CSR_valid)begin
        #10;
    end
    #26000;
    if(PE_pixels_0_0!==16'hffd0) $display("ERROR! at (0,0)\n");
if(PE_pixels_1_0!==16'h0048) $display("ERROR! at (1,0)\n");
if(PE_pixels_2_0!==16'h0018) $display("ERROR! at (2,0)\n");
if(PE_pixels_3_0!==16'h00e8) $display("ERROR! at (3,0)\n");
if(PE_pixels_4_0!==16'h001c) $display("ERROR! at (4,0)\n");
if(PE_pixels_5_0!==16'h001c) $display("ERROR! at (5,0)\n");
if(PE_pixels_6_0!==16'hff54) $display("ERROR! at (6,0)\n");
if(PE_pixels_7_0!==16'hfea4) $display("ERROR! at (7,0)\n");
if(PE_pixels_8_0!==16'hfda4) $display("ERROR! at (8,0)\n");
if(PE_pixels_9_0!==16'h0070) $display("ERROR! at (9,0)\n");
if(PE_pixels_10_0!==16'hff8c) $display("ERROR! at (10,0)\n");
if(PE_pixels_11_0!==16'hffd8) $display("ERROR! at (11,0)\n");
if(PE_pixels_12_0!==16'hffd0) $display("ERROR! at (12,0)\n");
if(PE_pixels_13_0!==16'hfe60) $display("ERROR! at (13,0)\n");
if(PE_pixels_14_0!==16'h012c) $display("ERROR! at (14,0)\n");
if(PE_pixels_15_0!==16'hfee2) $display("ERROR! at (15,0)\n");
if(PE_pixels_16_0!==16'hffe2) $display("ERROR! at (16,0)\n");
if(PE_pixels_17_0!==16'hfbd6) $display("ERROR! at (17,0)\n");
if(PE_pixels_18_0!==16'h00e6) $display("ERROR! at (18,0)\n");
if(PE_pixels_19_0!==16'h00f4) $display("ERROR! at (19,0)\n");
if(PE_pixels_20_0!==16'h01f8) $display("ERROR! at (20,0)\n");
if(PE_pixels_21_0!==16'h01b8) $display("ERROR! at (21,0)\n");
if(PE_pixels_22_0!==16'hffec) $display("ERROR! at (22,0)\n");
if(PE_pixels_23_0!==16'hffea) $display("ERROR! at (23,0)\n");
if(PE_pixels_24_0!==16'hfffe) $display("ERROR! at (24,0)\n");
if(PE_pixels_25_0!==16'hffec) $display("ERROR! at (25,0)\n");
if(PE_pixels_26_0!==16'h0004) $display("ERROR! at (26,0)\n");
if(PE_pixels_27_0!==16'h0000) $display("ERROR! at (27,0)\n");
if(PE_pixels_28_0!==16'h0000) $display("ERROR! at (28,0)\n");
if(PE_pixels_29_0!==16'h0000) $display("ERROR! at (29,0)\n");
if(PE_pixels_30_0!==16'h0000) $display("ERROR! at (30,0)\n");
if(PE_pixels_31_0!==16'h0000) $display("ERROR! at (31,0)\n");
if(PE_pixels_0_1!==16'hff70) $display("ERROR! at (0,1)\n");
if(PE_pixels_1_1!==16'h0034) $display("ERROR! at (1,1)\n");
if(PE_pixels_2_1!==16'h0084) $display("ERROR! at (2,1)\n");
if(PE_pixels_3_1!==16'hff6c) $display("ERROR! at (3,1)\n");
if(PE_pixels_4_1!==16'h0266) $display("ERROR! at (4,1)\n");
if(PE_pixels_5_1!==16'h014a) $display("ERROR! at (5,1)\n");
if(PE_pixels_6_1!==16'hfe00) $display("ERROR! at (6,1)\n");
if(PE_pixels_7_1!==16'hfc8e) $display("ERROR! at (7,1)\n");
if(PE_pixels_8_1!==16'hfc4e) $display("ERROR! at (8,1)\n");
if(PE_pixels_9_1!==16'hfb78) $display("ERROR! at (9,1)\n");
if(PE_pixels_10_1!==16'h0098) $display("ERROR! at (10,1)\n");
if(PE_pixels_11_1!==16'hfe12) $display("ERROR! at (11,1)\n");
if(PE_pixels_12_1!==16'hfdc6) $display("ERROR! at (12,1)\n");
if(PE_pixels_13_1!==16'hff20) $display("ERROR! at (13,1)\n");
if(PE_pixels_14_1!==16'h004c) $display("ERROR! at (14,1)\n");
if(PE_pixels_15_1!==16'hfe79) $display("ERROR! at (15,1)\n");
if(PE_pixels_16_1!==16'hfc54) $display("ERROR! at (16,1)\n");
if(PE_pixels_17_1!==16'hfdd9) $display("ERROR! at (17,1)\n");
if(PE_pixels_18_1!==16'hfacb) $display("ERROR! at (18,1)\n");
if(PE_pixels_19_1!==16'h0306) $display("ERROR! at (19,1)\n");
if(PE_pixels_20_1!==16'h03f9) $display("ERROR! at (20,1)\n");
if(PE_pixels_21_1!==16'h04d6) $display("ERROR! at (21,1)\n");
if(PE_pixels_22_1!==16'h0716) $display("ERROR! at (22,1)\n");
if(PE_pixels_23_1!==16'h0005) $display("ERROR! at (23,1)\n");
if(PE_pixels_24_1!==16'hffb2) $display("ERROR! at (24,1)\n");
if(PE_pixels_25_1!==16'hffe8) $display("ERROR! at (25,1)\n");
if(PE_pixels_26_1!==16'hff09) $display("ERROR! at (26,1)\n");
if(PE_pixels_27_1!==16'h0024) $display("ERROR! at (27,1)\n");
if(PE_pixels_28_1!==16'hffd8) $display("ERROR! at (28,1)\n");
if(PE_pixels_29_1!==16'h0008) $display("ERROR! at (29,1)\n");
if(PE_pixels_30_1!==16'h0000) $display("ERROR! at (30,1)\n");
if(PE_pixels_31_1!==16'h0000) $display("ERROR! at (31,1)\n");
if(PE_pixels_0_2!==16'h0050) $display("ERROR! at (0,2)\n");
if(PE_pixels_1_2!==16'hffd0) $display("ERROR! at (1,2)\n");
if(PE_pixels_2_2!==16'hfe66) $display("ERROR! at (2,2)\n");
if(PE_pixels_3_2!==16'h0034) $display("ERROR! at (3,2)\n");
if(PE_pixels_4_2!==16'hff60) $display("ERROR! at (4,2)\n");
if(PE_pixels_5_2!==16'h0065) $display("ERROR! at (5,2)\n");
if(PE_pixels_6_2!==16'h0116) $display("ERROR! at (6,2)\n");
if(PE_pixels_7_2!==16'hfec4) $display("ERROR! at (7,2)\n");
if(PE_pixels_8_2!==16'hf88b) $display("ERROR! at (8,2)\n");
if(PE_pixels_9_2!==16'hfe78) $display("ERROR! at (9,2)\n");
if(PE_pixels_10_2!==16'hffc8) $display("ERROR! at (10,2)\n");
if(PE_pixels_11_2!==16'h016a) $display("ERROR! at (11,2)\n");
if(PE_pixels_12_2!==16'hffd0) $display("ERROR! at (12,2)\n");
if(PE_pixels_13_2!==16'hfd0c) $display("ERROR! at (13,2)\n");
if(PE_pixels_14_2!==16'hff3e) $display("ERROR! at (14,2)\n");
if(PE_pixels_15_2!==16'h011e) $display("ERROR! at (15,2)\n");
if(PE_pixels_16_2!==16'h0033) $display("ERROR! at (16,2)\n");
if(PE_pixels_17_2!==16'hfe84) $display("ERROR! at (17,2)\n");
if(PE_pixels_18_2!==16'hfd44) $display("ERROR! at (18,2)\n");
if(PE_pixels_19_2!==16'h015e) $display("ERROR! at (19,2)\n");
if(PE_pixels_20_2!==16'h04fd) $display("ERROR! at (20,2)\n");
if(PE_pixels_21_2!==16'h078e) $display("ERROR! at (21,2)\n");
if(PE_pixels_22_2!==16'h04dc) $display("ERROR! at (22,2)\n");
if(PE_pixels_23_2!==16'h0794) $display("ERROR! at (23,2)\n");
if(PE_pixels_24_2!==16'hffd8) $display("ERROR! at (24,2)\n");
if(PE_pixels_25_2!==16'hff43) $display("ERROR! at (25,2)\n");
if(PE_pixels_26_2!==16'h007e) $display("ERROR! at (26,2)\n");
if(PE_pixels_27_2!==16'hfd76) $display("ERROR! at (27,2)\n");
if(PE_pixels_28_2!==16'hff54) $display("ERROR! at (28,2)\n");
if(PE_pixels_29_2!==16'hfd62) $display("ERROR! at (29,2)\n");
if(PE_pixels_30_2!==16'hfee0) $display("ERROR! at (30,2)\n");
if(PE_pixels_31_2!==16'h0050) $display("ERROR! at (31,2)\n");
if(PE_pixels_0_3!==16'h0074) $display("ERROR! at (0,3)\n");
if(PE_pixels_1_3!==16'h01da) $display("ERROR! at (1,3)\n");
if(PE_pixels_2_3!==16'h01c8) $display("ERROR! at (2,3)\n");
if(PE_pixels_3_3!==16'hfe0e) $display("ERROR! at (3,3)\n");
if(PE_pixels_4_3!==16'hfffa) $display("ERROR! at (4,3)\n");
if(PE_pixels_5_3!==16'h008c) $display("ERROR! at (5,3)\n");
if(PE_pixels_6_3!==16'hff9f) $display("ERROR! at (6,3)\n");
if(PE_pixels_7_3!==16'hfd4a) $display("ERROR! at (7,3)\n");
if(PE_pixels_8_3!==16'hfe02) $display("ERROR! at (8,3)\n");
if(PE_pixels_9_3!==16'hf9eb) $display("ERROR! at (9,3)\n");
if(PE_pixels_10_3!==16'h0061) $display("ERROR! at (10,3)\n");
if(PE_pixels_11_3!==16'h00aa) $display("ERROR! at (11,3)\n");
if(PE_pixels_12_3!==16'h009e) $display("ERROR! at (12,3)\n");
if(PE_pixels_13_3!==16'h0273) $display("ERROR! at (13,3)\n");
if(PE_pixels_14_3!==16'hf945) $display("ERROR! at (14,3)\n");
if(PE_pixels_15_3!==16'hfff0) $display("ERROR! at (15,3)\n");
if(PE_pixels_16_3!==16'hf958) $display("ERROR! at (16,3)\n");
if(PE_pixels_17_3!==16'h0700) $display("ERROR! at (17,3)\n");
if(PE_pixels_18_3!==16'hfec6) $display("ERROR! at (18,3)\n");
if(PE_pixels_19_3!==16'h0392) $display("ERROR! at (19,3)\n");
if(PE_pixels_20_3!==16'hfda6) $display("ERROR! at (20,3)\n");
if(PE_pixels_21_3!==16'hfecd) $display("ERROR! at (21,3)\n");
if(PE_pixels_22_3!==16'h06ae) $display("ERROR! at (22,3)\n");
if(PE_pixels_23_3!==16'h064b) $display("ERROR! at (23,3)\n");
if(PE_pixels_24_3!==16'h0366) $display("ERROR! at (24,3)\n");
if(PE_pixels_25_3!==16'h04a9) $display("ERROR! at (25,3)\n");
if(PE_pixels_26_3!==16'h00b7) $display("ERROR! at (26,3)\n");
if(PE_pixels_27_3!==16'h00e3) $display("ERROR! at (27,3)\n");
if(PE_pixels_28_3!==16'hfdcd) $display("ERROR! at (28,3)\n");
if(PE_pixels_29_3!==16'hfcdc) $display("ERROR! at (29,3)\n");
if(PE_pixels_30_3!==16'hfb3c) $display("ERROR! at (30,3)\n");
if(PE_pixels_31_3!==16'hfd44) $display("ERROR! at (31,3)\n");
if(PE_pixels_0_4!==16'hfeec) $display("ERROR! at (0,4)\n");
if(PE_pixels_1_4!==16'hfe7a) $display("ERROR! at (1,4)\n");
if(PE_pixels_2_4!==16'hfde4) $display("ERROR! at (2,4)\n");
if(PE_pixels_3_4!==16'h02a0) $display("ERROR! at (3,4)\n");
if(PE_pixels_4_4!==16'h00dd) $display("ERROR! at (4,4)\n");
if(PE_pixels_5_4!==16'h0124) $display("ERROR! at (5,4)\n");
if(PE_pixels_6_4!==16'h057f) $display("ERROR! at (6,4)\n");
if(PE_pixels_7_4!==16'h0666) $display("ERROR! at (7,4)\n");
if(PE_pixels_8_4!==16'hfc78) $display("ERROR! at (8,4)\n");
if(PE_pixels_9_4!==16'hf802) $display("ERROR! at (9,4)\n");
if(PE_pixels_10_4!==16'hff1e) $display("ERROR! at (10,4)\n");
if(PE_pixels_11_4!==16'h01ce) $display("ERROR! at (11,4)\n");
if(PE_pixels_12_4!==16'h042b) $display("ERROR! at (12,4)\n");
if(PE_pixels_13_4!==16'hfcfa) $display("ERROR! at (13,4)\n");
if(PE_pixels_14_4!==16'hfcc2) $display("ERROR! at (14,4)\n");
if(PE_pixels_15_4!==16'hff83) $display("ERROR! at (15,4)\n");
if(PE_pixels_16_4!==16'h0525) $display("ERROR! at (16,4)\n");
if(PE_pixels_17_4!==16'h020a) $display("ERROR! at (17,4)\n");
if(PE_pixels_18_4!==16'hf744) $display("ERROR! at (18,4)\n");
if(PE_pixels_19_4!==16'hfc98) $display("ERROR! at (19,4)\n");
if(PE_pixels_20_4!==16'hfd4e) $display("ERROR! at (20,4)\n");
if(PE_pixels_21_4!==16'hff2d) $display("ERROR! at (21,4)\n");
if(PE_pixels_22_4!==16'hf971) $display("ERROR! at (22,4)\n");
if(PE_pixels_23_4!==16'h0629) $display("ERROR! at (23,4)\n");
if(PE_pixels_24_4!==16'h03d5) $display("ERROR! at (24,4)\n");
if(PE_pixels_25_4!==16'h003c) $display("ERROR! at (25,4)\n");
if(PE_pixels_26_4!==16'h0a4a) $display("ERROR! at (26,4)\n");
if(PE_pixels_27_4!==16'h02f9) $display("ERROR! at (27,4)\n");
if(PE_pixels_28_4!==16'h02f2) $display("ERROR! at (28,4)\n");
if(PE_pixels_29_4!==16'h0110) $display("ERROR! at (29,4)\n");
if(PE_pixels_30_4!==16'hfcb4) $display("ERROR! at (30,4)\n");
if(PE_pixels_31_4!==16'hfe98) $display("ERROR! at (31,4)\n");
if(PE_pixels_0_5!==16'h00a6) $display("ERROR! at (0,5)\n");
if(PE_pixels_1_5!==16'h0092) $display("ERROR! at (1,5)\n");
if(PE_pixels_2_5!==16'h00ec) $display("ERROR! at (2,5)\n");
if(PE_pixels_3_5!==16'hfd7a) $display("ERROR! at (3,5)\n");
if(PE_pixels_4_5!==16'h00eb) $display("ERROR! at (4,5)\n");
if(PE_pixels_5_5!==16'hfd17) $display("ERROR! at (5,5)\n");
if(PE_pixels_6_5!==16'h0154) $display("ERROR! at (6,5)\n");
if(PE_pixels_7_5!==16'hfbeb) $display("ERROR! at (7,5)\n");
if(PE_pixels_8_5!==16'h04a8) $display("ERROR! at (8,5)\n");
if(PE_pixels_9_5!==16'h0129) $display("ERROR! at (9,5)\n");
if(PE_pixels_10_5!==16'h01f3) $display("ERROR! at (10,5)\n");
if(PE_pixels_11_5!==16'hffa3) $display("ERROR! at (11,5)\n");
if(PE_pixels_12_5!==16'h026c) $display("ERROR! at (12,5)\n");
if(PE_pixels_13_5!==16'hff46) $display("ERROR! at (13,5)\n");
if(PE_pixels_14_5!==16'hfdd8) $display("ERROR! at (14,5)\n");
if(PE_pixels_15_5!==16'hfcf5) $display("ERROR! at (15,5)\n");
if(PE_pixels_16_5!==16'h00e0) $display("ERROR! at (16,5)\n");
if(PE_pixels_17_5!==16'h002b) $display("ERROR! at (17,5)\n");
if(PE_pixels_18_5!==16'h014c) $display("ERROR! at (18,5)\n");
if(PE_pixels_19_5!==16'h00e0) $display("ERROR! at (19,5)\n");
if(PE_pixels_20_5!==16'hfe08) $display("ERROR! at (20,5)\n");
if(PE_pixels_21_5!==16'hf8b0) $display("ERROR! at (21,5)\n");
if(PE_pixels_22_5!==16'hfdcf) $display("ERROR! at (22,5)\n");
if(PE_pixels_23_5!==16'hff5a) $display("ERROR! at (23,5)\n");
if(PE_pixels_24_5!==16'h0141) $display("ERROR! at (24,5)\n");
if(PE_pixels_25_5!==16'h0342) $display("ERROR! at (25,5)\n");
if(PE_pixels_26_5!==16'hfee8) $display("ERROR! at (26,5)\n");
if(PE_pixels_27_5!==16'hff51) $display("ERROR! at (27,5)\n");
if(PE_pixels_28_5!==16'hff8d) $display("ERROR! at (28,5)\n");
if(PE_pixels_29_5!==16'h04b6) $display("ERROR! at (29,5)\n");
if(PE_pixels_30_5!==16'h00d4) $display("ERROR! at (30,5)\n");
if(PE_pixels_31_5!==16'hfe5c) $display("ERROR! at (31,5)\n");
if(PE_pixels_0_6!==16'hff3a) $display("ERROR! at (0,6)\n");
if(PE_pixels_1_6!==16'h00aa) $display("ERROR! at (1,6)\n");
if(PE_pixels_2_6!==16'h01e0) $display("ERROR! at (2,6)\n");
if(PE_pixels_3_6!==16'h031a) $display("ERROR! at (3,6)\n");
if(PE_pixels_4_6!==16'h0318) $display("ERROR! at (4,6)\n");
if(PE_pixels_5_6!==16'hfb2f) $display("ERROR! at (5,6)\n");
if(PE_pixels_6_6!==16'h005d) $display("ERROR! at (6,6)\n");
if(PE_pixels_7_6!==16'hfebb) $display("ERROR! at (7,6)\n");
if(PE_pixels_8_6!==16'hfe6c) $display("ERROR! at (8,6)\n");
if(PE_pixels_9_6!==16'h0049) $display("ERROR! at (9,6)\n");
if(PE_pixels_10_6!==16'hffeb) $display("ERROR! at (10,6)\n");
if(PE_pixels_11_6!==16'h0218) $display("ERROR! at (11,6)\n");
if(PE_pixels_12_6!==16'h0145) $display("ERROR! at (12,6)\n");
if(PE_pixels_13_6!==16'hff50) $display("ERROR! at (13,6)\n");
if(PE_pixels_14_6!==16'h03e6) $display("ERROR! at (14,6)\n");
if(PE_pixels_15_6!==16'hfe8a) $display("ERROR! at (15,6)\n");
if(PE_pixels_16_6!==16'hff4c) $display("ERROR! at (16,6)\n");
if(PE_pixels_17_6!==16'hfe60) $display("ERROR! at (17,6)\n");
if(PE_pixels_18_6!==16'hffe9) $display("ERROR! at (18,6)\n");
if(PE_pixels_19_6!==16'hfdb8) $display("ERROR! at (19,6)\n");
if(PE_pixels_20_6!==16'h0252) $display("ERROR! at (20,6)\n");
if(PE_pixels_21_6!==16'hf694) $display("ERROR! at (21,6)\n");
if(PE_pixels_22_6!==16'h04be) $display("ERROR! at (22,6)\n");
if(PE_pixels_23_6!==16'h0205) $display("ERROR! at (23,6)\n");
if(PE_pixels_24_6!==16'h04b6) $display("ERROR! at (24,6)\n");
if(PE_pixels_25_6!==16'hfb65) $display("ERROR! at (25,6)\n");
if(PE_pixels_26_6!==16'h04c4) $display("ERROR! at (26,6)\n");
if(PE_pixels_27_6!==16'h0210) $display("ERROR! at (27,6)\n");
if(PE_pixels_28_6!==16'hfee7) $display("ERROR! at (28,6)\n");
if(PE_pixels_29_6!==16'h011a) $display("ERROR! at (29,6)\n");
if(PE_pixels_30_6!==16'hfe88) $display("ERROR! at (30,6)\n");
if(PE_pixels_31_6!==16'hfe84) $display("ERROR! at (31,6)\n");
if(PE_pixels_0_7!==16'hfdf8) $display("ERROR! at (0,7)\n");
if(PE_pixels_1_7!==16'hff9d) $display("ERROR! at (1,7)\n");
if(PE_pixels_2_7!==16'h024c) $display("ERROR! at (2,7)\n");
if(PE_pixels_3_7!==16'h010c) $display("ERROR! at (3,7)\n");
if(PE_pixels_4_7!==16'h0806) $display("ERROR! at (4,7)\n");
if(PE_pixels_5_7!==16'h0313) $display("ERROR! at (5,7)\n");
if(PE_pixels_6_7!==16'h0172) $display("ERROR! at (6,7)\n");
if(PE_pixels_7_7!==16'h0002) $display("ERROR! at (7,7)\n");
if(PE_pixels_8_7!==16'hfbe5) $display("ERROR! at (8,7)\n");
if(PE_pixels_9_7!==16'h0002) $display("ERROR! at (9,7)\n");
if(PE_pixels_10_7!==16'h0093) $display("ERROR! at (10,7)\n");
if(PE_pixels_11_7!==16'h0595) $display("ERROR! at (11,7)\n");
if(PE_pixels_12_7!==16'hff4f) $display("ERROR! at (12,7)\n");
if(PE_pixels_13_7!==16'h00ad) $display("ERROR! at (13,7)\n");
if(PE_pixels_14_7!==16'h033e) $display("ERROR! at (14,7)\n");
if(PE_pixels_15_7!==16'h0000) $display("ERROR! at (15,7)\n");
if(PE_pixels_16_7!==16'h0360) $display("ERROR! at (16,7)\n");
if(PE_pixels_17_7!==16'h00f3) $display("ERROR! at (17,7)\n");
if(PE_pixels_18_7!==16'hfdfe) $display("ERROR! at (18,7)\n");
if(PE_pixels_19_7!==16'h009b) $display("ERROR! at (19,7)\n");
if(PE_pixels_20_7!==16'h017b) $display("ERROR! at (20,7)\n");
if(PE_pixels_21_7!==16'hfd69) $display("ERROR! at (21,7)\n");
if(PE_pixels_22_7!==16'hff34) $display("ERROR! at (22,7)\n");
if(PE_pixels_23_7!==16'hfc8f) $display("ERROR! at (23,7)\n");
if(PE_pixels_24_7!==16'hfffc) $display("ERROR! at (24,7)\n");
if(PE_pixels_25_7!==16'hfef5) $display("ERROR! at (25,7)\n");
if(PE_pixels_26_7!==16'h08a4) $display("ERROR! at (26,7)\n");
if(PE_pixels_27_7!==16'hfbd4) $display("ERROR! at (27,7)\n");
if(PE_pixels_28_7!==16'hfe10) $display("ERROR! at (28,7)\n");
if(PE_pixels_29_7!==16'hfd7a) $display("ERROR! at (29,7)\n");
if(PE_pixels_30_7!==16'hfd44) $display("ERROR! at (30,7)\n");
if(PE_pixels_31_7!==16'h0000) $display("ERROR! at (31,7)\n");
if(PE_pixels_0_8!==16'hff32) $display("ERROR! at (0,8)\n");
if(PE_pixels_1_8!==16'hfc86) $display("ERROR! at (1,8)\n");
if(PE_pixels_2_8!==16'hff6d) $display("ERROR! at (2,8)\n");
if(PE_pixels_3_8!==16'h05de) $display("ERROR! at (3,8)\n");
if(PE_pixels_4_8!==16'h032f) $display("ERROR! at (4,8)\n");
if(PE_pixels_5_8!==16'h033d) $display("ERROR! at (5,8)\n");
if(PE_pixels_6_8!==16'h020c) $display("ERROR! at (6,8)\n");
if(PE_pixels_7_8!==16'h0705) $display("ERROR! at (7,8)\n");
if(PE_pixels_8_8!==16'hfb9e) $display("ERROR! at (8,8)\n");
if(PE_pixels_9_8!==16'hffd0) $display("ERROR! at (9,8)\n");
if(PE_pixels_10_8!==16'hfd3b) $display("ERROR! at (10,8)\n");
if(PE_pixels_11_8!==16'hff7c) $display("ERROR! at (11,8)\n");
if(PE_pixels_12_8!==16'h01d6) $display("ERROR! at (12,8)\n");
if(PE_pixels_13_8!==16'hff89) $display("ERROR! at (13,8)\n");
if(PE_pixels_14_8!==16'hfe8b) $display("ERROR! at (14,8)\n");
if(PE_pixels_15_8!==16'hff1e) $display("ERROR! at (15,8)\n");
if(PE_pixels_16_8!==16'h008c) $display("ERROR! at (16,8)\n");
if(PE_pixels_17_8!==16'hfd6b) $display("ERROR! at (17,8)\n");
if(PE_pixels_18_8!==16'h03a4) $display("ERROR! at (18,8)\n");
if(PE_pixels_19_8!==16'hfeb9) $display("ERROR! at (19,8)\n");
if(PE_pixels_20_8!==16'h0422) $display("ERROR! at (20,8)\n");
if(PE_pixels_21_8!==16'hfa50) $display("ERROR! at (21,8)\n");
if(PE_pixels_22_8!==16'h0148) $display("ERROR! at (22,8)\n");
if(PE_pixels_23_8!==16'hfe0f) $display("ERROR! at (23,8)\n");
if(PE_pixels_24_8!==16'hfe88) $display("ERROR! at (24,8)\n");
if(PE_pixels_25_8!==16'h03d6) $display("ERROR! at (25,8)\n");
if(PE_pixels_26_8!==16'h0117) $display("ERROR! at (26,8)\n");
if(PE_pixels_27_8!==16'h046f) $display("ERROR! at (27,8)\n");
if(PE_pixels_28_8!==16'hfbd3) $display("ERROR! at (28,8)\n");
if(PE_pixels_29_8!==16'hfcb4) $display("ERROR! at (29,8)\n");
if(PE_pixels_30_8!==16'hf81b) $display("ERROR! at (30,8)\n");
if(PE_pixels_31_8!==16'h0048) $display("ERROR! at (31,8)\n");
if(PE_pixels_0_9!==16'h00ab) $display("ERROR! at (0,9)\n");
if(PE_pixels_1_9!==16'hfee8) $display("ERROR! at (1,9)\n");
if(PE_pixels_2_9!==16'h00c4) $display("ERROR! at (2,9)\n");
if(PE_pixels_3_9!==16'hfb9f) $display("ERROR! at (3,9)\n");
if(PE_pixels_4_9!==16'h08af) $display("ERROR! at (4,9)\n");
if(PE_pixels_5_9!==16'h07e9) $display("ERROR! at (5,9)\n");
if(PE_pixels_6_9!==16'h022a) $display("ERROR! at (6,9)\n");
if(PE_pixels_7_9!==16'h018a) $display("ERROR! at (7,9)\n");
if(PE_pixels_8_9!==16'hff5a) $display("ERROR! at (8,9)\n");
if(PE_pixels_9_9!==16'hfab8) $display("ERROR! at (9,9)\n");
if(PE_pixels_10_9!==16'hfd24) $display("ERROR! at (10,9)\n");
if(PE_pixels_11_9!==16'hff60) $display("ERROR! at (11,9)\n");
if(PE_pixels_12_9!==16'hfe35) $display("ERROR! at (12,9)\n");
if(PE_pixels_13_9!==16'h005b) $display("ERROR! at (13,9)\n");
if(PE_pixels_14_9!==16'h0139) $display("ERROR! at (14,9)\n");
if(PE_pixels_15_9!==16'hfed3) $display("ERROR! at (15,9)\n");
if(PE_pixels_16_9!==16'hffcd) $display("ERROR! at (16,9)\n");
if(PE_pixels_17_9!==16'h02c2) $display("ERROR! at (17,9)\n");
if(PE_pixels_18_9!==16'hff6c) $display("ERROR! at (18,9)\n");
if(PE_pixels_19_9!==16'hfe88) $display("ERROR! at (19,9)\n");
if(PE_pixels_20_9!==16'hfe12) $display("ERROR! at (20,9)\n");
if(PE_pixels_21_9!==16'hfc4a) $display("ERROR! at (21,9)\n");
if(PE_pixels_22_9!==16'hfd6c) $display("ERROR! at (22,9)\n");
if(PE_pixels_23_9!==16'hfffd) $display("ERROR! at (23,9)\n");
if(PE_pixels_24_9!==16'h001f) $display("ERROR! at (24,9)\n");
if(PE_pixels_25_9!==16'hff8e) $display("ERROR! at (25,9)\n");
if(PE_pixels_26_9!==16'h0343) $display("ERROR! at (26,9)\n");
if(PE_pixels_27_9!==16'h049a) $display("ERROR! at (27,9)\n");
if(PE_pixels_28_9!==16'hfe86) $display("ERROR! at (28,9)\n");
if(PE_pixels_29_9!==16'hff8d) $display("ERROR! at (29,9)\n");
if(PE_pixels_30_9!==16'hfaad) $display("ERROR! at (30,9)\n");
if(PE_pixels_31_9!==16'hfd9a) $display("ERROR! at (31,9)\n");
if(PE_pixels_0_10!==16'hff5d) $display("ERROR! at (0,10)\n");
if(PE_pixels_1_10!==16'hfd95) $display("ERROR! at (1,10)\n");
if(PE_pixels_2_10!==16'hfd36) $display("ERROR! at (2,10)\n");
if(PE_pixels_3_10!==16'h0450) $display("ERROR! at (3,10)\n");
if(PE_pixels_4_10!==16'h03a7) $display("ERROR! at (4,10)\n");
if(PE_pixels_5_10!==16'h0318) $display("ERROR! at (5,10)\n");
if(PE_pixels_6_10!==16'h059f) $display("ERROR! at (6,10)\n");
if(PE_pixels_7_10!==16'h00ac) $display("ERROR! at (7,10)\n");
if(PE_pixels_8_10!==16'h024f) $display("ERROR! at (8,10)\n");
if(PE_pixels_9_10!==16'h0061) $display("ERROR! at (9,10)\n");
if(PE_pixels_10_10!==16'h0435) $display("ERROR! at (10,10)\n");
if(PE_pixels_11_10!==16'hf959) $display("ERROR! at (11,10)\n");
if(PE_pixels_12_10!==16'hfd3e) $display("ERROR! at (12,10)\n");
if(PE_pixels_13_10!==16'hff99) $display("ERROR! at (13,10)\n");
if(PE_pixels_14_10!==16'hfea7) $display("ERROR! at (14,10)\n");
if(PE_pixels_15_10!==16'hfeed) $display("ERROR! at (15,10)\n");
if(PE_pixels_16_10!==16'h015c) $display("ERROR! at (16,10)\n");
if(PE_pixels_17_10!==16'h006d) $display("ERROR! at (17,10)\n");
if(PE_pixels_18_10!==16'h046d) $display("ERROR! at (18,10)\n");
if(PE_pixels_19_10!==16'hfd68) $display("ERROR! at (19,10)\n");
if(PE_pixels_20_10!==16'h0029) $display("ERROR! at (20,10)\n");
if(PE_pixels_21_10!==16'hfd0a) $display("ERROR! at (21,10)\n");
if(PE_pixels_22_10!==16'hfc64) $display("ERROR! at (22,10)\n");
if(PE_pixels_23_10!==16'hfe97) $display("ERROR! at (23,10)\n");
if(PE_pixels_24_10!==16'hfb41) $display("ERROR! at (24,10)\n");
if(PE_pixels_25_10!==16'h0557) $display("ERROR! at (25,10)\n");
if(PE_pixels_26_10!==16'hf812) $display("ERROR! at (26,10)\n");
if(PE_pixels_27_10!==16'h08ec) $display("ERROR! at (27,10)\n");
if(PE_pixels_28_10!==16'hfed9) $display("ERROR! at (28,10)\n");
if(PE_pixels_29_10!==16'h05b7) $display("ERROR! at (29,10)\n");
if(PE_pixels_30_10!==16'hf8dd) $display("ERROR! at (30,10)\n");
if(PE_pixels_31_10!==16'hfe34) $display("ERROR! at (31,10)\n");
if(PE_pixels_0_11!==16'h0176) $display("ERROR! at (0,11)\n");
if(PE_pixels_1_11!==16'hff93) $display("ERROR! at (1,11)\n");
if(PE_pixels_2_11!==16'hfdb1) $display("ERROR! at (2,11)\n");
if(PE_pixels_3_11!==16'hf8c5) $display("ERROR! at (3,11)\n");
if(PE_pixels_4_11!==16'hfe90) $display("ERROR! at (4,11)\n");
if(PE_pixels_5_11!==16'h0880) $display("ERROR! at (5,11)\n");
if(PE_pixels_6_11!==16'h03e2) $display("ERROR! at (6,11)\n");
if(PE_pixels_7_11!==16'h026f) $display("ERROR! at (7,11)\n");
if(PE_pixels_8_11!==16'h0242) $display("ERROR! at (8,11)\n");
if(PE_pixels_9_11!==16'h01e3) $display("ERROR! at (9,11)\n");
if(PE_pixels_10_11!==16'hfddb) $display("ERROR! at (10,11)\n");
if(PE_pixels_11_11!==16'h011b) $display("ERROR! at (11,11)\n");
if(PE_pixels_12_11!==16'hfd01) $display("ERROR! at (12,11)\n");
if(PE_pixels_13_11!==16'hfe8b) $display("ERROR! at (13,11)\n");
if(PE_pixels_14_11!==16'h0046) $display("ERROR! at (14,11)\n");
if(PE_pixels_15_11!==16'hff5b) $display("ERROR! at (15,11)\n");
if(PE_pixels_16_11!==16'h0718) $display("ERROR! at (16,11)\n");
if(PE_pixels_17_11!==16'h03df) $display("ERROR! at (17,11)\n");
if(PE_pixels_18_11!==16'hff00) $display("ERROR! at (18,11)\n");
if(PE_pixels_19_11!==16'h02db) $display("ERROR! at (19,11)\n");
if(PE_pixels_20_11!==16'h019f) $display("ERROR! at (20,11)\n");
if(PE_pixels_21_11!==16'h02c3) $display("ERROR! at (21,11)\n");
if(PE_pixels_22_11!==16'hfe55) $display("ERROR! at (22,11)\n");
if(PE_pixels_23_11!==16'h000f) $display("ERROR! at (23,11)\n");
if(PE_pixels_24_11!==16'hfc3f) $display("ERROR! at (24,11)\n");
if(PE_pixels_25_11!==16'hfbfd) $display("ERROR! at (25,11)\n");
if(PE_pixels_26_11!==16'h0231) $display("ERROR! at (26,11)\n");
if(PE_pixels_27_11!==16'h0151) $display("ERROR! at (27,11)\n");
if(PE_pixels_28_11!==16'h060f) $display("ERROR! at (28,11)\n");
if(PE_pixels_29_11!==16'hff13) $display("ERROR! at (29,11)\n");
if(PE_pixels_30_11!==16'hff6c) $display("ERROR! at (30,11)\n");
if(PE_pixels_31_11!==16'hfe1b) $display("ERROR! at (31,11)\n");
if(PE_pixels_0_12!==16'h002e) $display("ERROR! at (0,12)\n");
if(PE_pixels_1_12!==16'hfe8a) $display("ERROR! at (1,12)\n");
if(PE_pixels_2_12!==16'h000e) $display("ERROR! at (2,12)\n");
if(PE_pixels_3_12!==16'hffc2) $display("ERROR! at (3,12)\n");
if(PE_pixels_4_12!==16'h0368) $display("ERROR! at (4,12)\n");
if(PE_pixels_5_12!==16'hffcc) $display("ERROR! at (5,12)\n");
if(PE_pixels_6_12!==16'h04bb) $display("ERROR! at (6,12)\n");
if(PE_pixels_7_12!==16'h0244) $display("ERROR! at (7,12)\n");
if(PE_pixels_8_12!==16'h018f) $display("ERROR! at (8,12)\n");
if(PE_pixels_9_12!==16'h0240) $display("ERROR! at (9,12)\n");
if(PE_pixels_10_12!==16'h00d8) $display("ERROR! at (10,12)\n");
if(PE_pixels_11_12!==16'h03d9) $display("ERROR! at (11,12)\n");
if(PE_pixels_12_12!==16'hfcff) $display("ERROR! at (12,12)\n");
if(PE_pixels_13_12!==16'hfb8e) $display("ERROR! at (13,12)\n");
if(PE_pixels_14_12!==16'h000a) $display("ERROR! at (14,12)\n");
if(PE_pixels_15_12!==16'h0234) $display("ERROR! at (15,12)\n");
if(PE_pixels_16_12!==16'h0072) $display("ERROR! at (16,12)\n");
if(PE_pixels_17_12!==16'h05fa) $display("ERROR! at (17,12)\n");
if(PE_pixels_18_12!==16'h07e3) $display("ERROR! at (18,12)\n");
if(PE_pixels_19_12!==16'hfe34) $display("ERROR! at (19,12)\n");
if(PE_pixels_20_12!==16'h004c) $display("ERROR! at (20,12)\n");
if(PE_pixels_21_12!==16'hfeb9) $display("ERROR! at (21,12)\n");
if(PE_pixels_22_12!==16'h0136) $display("ERROR! at (22,12)\n");
if(PE_pixels_23_12!==16'h0017) $display("ERROR! at (23,12)\n");
if(PE_pixels_24_12!==16'hfed7) $display("ERROR! at (24,12)\n");
if(PE_pixels_25_12!==16'hfdb8) $display("ERROR! at (25,12)\n");
if(PE_pixels_26_12!==16'hfcd8) $display("ERROR! at (26,12)\n");
if(PE_pixels_27_12!==16'hfffa) $display("ERROR! at (27,12)\n");
if(PE_pixels_28_12!==16'h0128) $display("ERROR! at (28,12)\n");
if(PE_pixels_29_12!==16'h0243) $display("ERROR! at (29,12)\n");
if(PE_pixels_30_12!==16'h0120) $display("ERROR! at (30,12)\n");
if(PE_pixels_31_12!==16'hfe14) $display("ERROR! at (31,12)\n");
if(PE_pixels_0_13!==16'h0110) $display("ERROR! at (0,13)\n");
if(PE_pixels_1_13!==16'hfdb5) $display("ERROR! at (1,13)\n");
if(PE_pixels_2_13!==16'hfdbc) $display("ERROR! at (2,13)\n");
if(PE_pixels_3_13!==16'hfda2) $display("ERROR! at (3,13)\n");
if(PE_pixels_4_13!==16'hfcbc) $display("ERROR! at (4,13)\n");
if(PE_pixels_5_13!==16'h07ec) $display("ERROR! at (5,13)\n");
if(PE_pixels_6_13!==16'h0404) $display("ERROR! at (6,13)\n");
if(PE_pixels_7_13!==16'h013d) $display("ERROR! at (7,13)\n");
if(PE_pixels_8_13!==16'h0273) $display("ERROR! at (8,13)\n");
if(PE_pixels_9_13!==16'hfd7b) $display("ERROR! at (9,13)\n");
if(PE_pixels_10_13!==16'h0207) $display("ERROR! at (10,13)\n");
if(PE_pixels_11_13!==16'h0196) $display("ERROR! at (11,13)\n");
if(PE_pixels_12_13!==16'h023f) $display("ERROR! at (12,13)\n");
if(PE_pixels_13_13!==16'hffb5) $display("ERROR! at (13,13)\n");
if(PE_pixels_14_13!==16'hfc35) $display("ERROR! at (14,13)\n");
if(PE_pixels_15_13!==16'hffef) $display("ERROR! at (15,13)\n");
if(PE_pixels_16_13!==16'h05fe) $display("ERROR! at (16,13)\n");
if(PE_pixels_17_13!==16'h068a) $display("ERROR! at (17,13)\n");
if(PE_pixels_18_13!==16'hff54) $display("ERROR! at (18,13)\n");
if(PE_pixels_19_13!==16'h00b8) $display("ERROR! at (19,13)\n");
if(PE_pixels_20_13!==16'hff1e) $display("ERROR! at (20,13)\n");
if(PE_pixels_21_13!==16'hffdb) $display("ERROR! at (21,13)\n");
if(PE_pixels_22_13!==16'hfeaa) $display("ERROR! at (22,13)\n");
if(PE_pixels_23_13!==16'hfff3) $display("ERROR! at (23,13)\n");
if(PE_pixels_24_13!==16'h00f9) $display("ERROR! at (24,13)\n");
if(PE_pixels_25_13!==16'hfed4) $display("ERROR! at (25,13)\n");
if(PE_pixels_26_13!==16'h0388) $display("ERROR! at (26,13)\n");
if(PE_pixels_27_13!==16'hf522) $display("ERROR! at (27,13)\n");
if(PE_pixels_28_13!==16'h039e) $display("ERROR! at (28,13)\n");
if(PE_pixels_29_13!==16'h031e) $display("ERROR! at (29,13)\n");
if(PE_pixels_30_13!==16'hffc4) $display("ERROR! at (30,13)\n");
if(PE_pixels_31_13!==16'h0143) $display("ERROR! at (31,13)\n");
if(PE_pixels_0_14!==16'h0036) $display("ERROR! at (0,14)\n");
if(PE_pixels_1_14!==16'h018c) $display("ERROR! at (1,14)\n");
if(PE_pixels_2_14!==16'hfebe) $display("ERROR! at (2,14)\n");
if(PE_pixels_3_14!==16'hff7d) $display("ERROR! at (3,14)\n");
if(PE_pixels_4_14!==16'hfdc2) $display("ERROR! at (4,14)\n");
if(PE_pixels_5_14!==16'h010f) $display("ERROR! at (5,14)\n");
if(PE_pixels_6_14!==16'hffd5) $display("ERROR! at (6,14)\n");
if(PE_pixels_7_14!==16'h008a) $display("ERROR! at (7,14)\n");
if(PE_pixels_8_14!==16'h04e2) $display("ERROR! at (8,14)\n");
if(PE_pixels_9_14!==16'hfc5e) $display("ERROR! at (9,14)\n");
if(PE_pixels_10_14!==16'hff24) $display("ERROR! at (10,14)\n");
if(PE_pixels_11_14!==16'hffd2) $display("ERROR! at (11,14)\n");
if(PE_pixels_12_14!==16'h04e9) $display("ERROR! at (12,14)\n");
if(PE_pixels_13_14!==16'h02f5) $display("ERROR! at (13,14)\n");
if(PE_pixels_14_14!==16'hfffd) $display("ERROR! at (14,14)\n");
if(PE_pixels_15_14!==16'hfddf) $display("ERROR! at (15,14)\n");
if(PE_pixels_16_14!==16'hf6d3) $display("ERROR! at (16,14)\n");
if(PE_pixels_17_14!==16'h00a6) $display("ERROR! at (17,14)\n");
if(PE_pixels_18_14!==16'h0990) $display("ERROR! at (18,14)\n");
if(PE_pixels_19_14!==16'h0540) $display("ERROR! at (19,14)\n");
if(PE_pixels_20_14!==16'h003a) $display("ERROR! at (20,14)\n");
if(PE_pixels_21_14!==16'h00ca) $display("ERROR! at (21,14)\n");
if(PE_pixels_22_14!==16'hff2b) $display("ERROR! at (22,14)\n");
if(PE_pixels_23_14!==16'hfff5) $display("ERROR! at (23,14)\n");
if(PE_pixels_24_14!==16'h0200) $display("ERROR! at (24,14)\n");
if(PE_pixels_25_14!==16'hfe43) $display("ERROR! at (25,14)\n");
if(PE_pixels_26_14!==16'hf983) $display("ERROR! at (26,14)\n");
if(PE_pixels_27_14!==16'hfc27) $display("ERROR! at (27,14)\n");
if(PE_pixels_28_14!==16'hfe1c) $display("ERROR! at (28,14)\n");
if(PE_pixels_29_14!==16'hffb2) $display("ERROR! at (29,14)\n");
if(PE_pixels_30_14!==16'h0421) $display("ERROR! at (30,14)\n");
if(PE_pixels_31_14!==16'h00e1) $display("ERROR! at (31,14)\n");
if(PE_pixels_0_15!==16'hfe1f) $display("ERROR! at (0,15)\n");
if(PE_pixels_1_15!==16'h0246) $display("ERROR! at (1,15)\n");
if(PE_pixels_2_15!==16'hfedc) $display("ERROR! at (2,15)\n");
if(PE_pixels_3_15!==16'h0632) $display("ERROR! at (3,15)\n");
if(PE_pixels_4_15!==16'hfbbe) $display("ERROR! at (4,15)\n");
if(PE_pixels_5_15!==16'hffee) $display("ERROR! at (5,15)\n");
if(PE_pixels_6_15!==16'hff2d) $display("ERROR! at (6,15)\n");
if(PE_pixels_7_15!==16'hf9ef) $display("ERROR! at (7,15)\n");
if(PE_pixels_8_15!==16'h0665) $display("ERROR! at (8,15)\n");
if(PE_pixels_9_15!==16'hfebb) $display("ERROR! at (9,15)\n");
if(PE_pixels_10_15!==16'h0363) $display("ERROR! at (10,15)\n");
if(PE_pixels_11_15!==16'hfe1d) $display("ERROR! at (11,15)\n");
if(PE_pixels_12_15!==16'h02f4) $display("ERROR! at (12,15)\n");
if(PE_pixels_13_15!==16'h0397) $display("ERROR! at (13,15)\n");
if(PE_pixels_14_15!==16'hfee6) $display("ERROR! at (14,15)\n");
if(PE_pixels_15_15!==16'hf8f9) $display("ERROR! at (15,15)\n");
if(PE_pixels_16_15!==16'hfec5) $display("ERROR! at (16,15)\n");
if(PE_pixels_17_15!==16'h0145) $display("ERROR! at (17,15)\n");
if(PE_pixels_18_15!==16'h0292) $display("ERROR! at (18,15)\n");
if(PE_pixels_19_15!==16'h0398) $display("ERROR! at (19,15)\n");
if(PE_pixels_20_15!==16'hffc7) $display("ERROR! at (20,15)\n");
if(PE_pixels_21_15!==16'h00e0) $display("ERROR! at (21,15)\n");
if(PE_pixels_22_15!==16'hfeae) $display("ERROR! at (22,15)\n");
if(PE_pixels_23_15!==16'hff46) $display("ERROR! at (23,15)\n");
if(PE_pixels_24_15!==16'h0207) $display("ERROR! at (24,15)\n");
if(PE_pixels_25_15!==16'hff6a) $display("ERROR! at (25,15)\n");
if(PE_pixels_26_15!==16'h00d7) $display("ERROR! at (26,15)\n");
if(PE_pixels_27_15!==16'hfade) $display("ERROR! at (27,15)\n");
if(PE_pixels_28_15!==16'hf70b) $display("ERROR! at (28,15)\n");
if(PE_pixels_29_15!==16'h00da) $display("ERROR! at (29,15)\n");
if(PE_pixels_30_15!==16'hfce4) $display("ERROR! at (30,15)\n");
if(PE_pixels_31_15!==16'h0007) $display("ERROR! at (31,15)\n");
if(PE_pixels_0_16!==16'hfff5) $display("ERROR! at (0,16)\n");
if(PE_pixels_1_16!==16'hff72) $display("ERROR! at (1,16)\n");
if(PE_pixels_2_16!==16'hff0f) $display("ERROR! at (2,16)\n");
if(PE_pixels_3_16!==16'hfdb6) $display("ERROR! at (3,16)\n");
if(PE_pixels_4_16!==16'h01ba) $display("ERROR! at (4,16)\n");
if(PE_pixels_5_16!==16'h0324) $display("ERROR! at (5,16)\n");
if(PE_pixels_6_16!==16'hff4e) $display("ERROR! at (6,16)\n");
if(PE_pixels_7_16!==16'hfe2a) $display("ERROR! at (7,16)\n");
if(PE_pixels_8_16!==16'h02b4) $display("ERROR! at (8,16)\n");
if(PE_pixels_9_16!==16'hfde8) $display("ERROR! at (9,16)\n");
if(PE_pixels_10_16!==16'hfe86) $display("ERROR! at (10,16)\n");
if(PE_pixels_11_16!==16'hfd9b) $display("ERROR! at (11,16)\n");
if(PE_pixels_12_16!==16'h0427) $display("ERROR! at (12,16)\n");
if(PE_pixels_13_16!==16'h07ec) $display("ERROR! at (13,16)\n");
if(PE_pixels_14_16!==16'hfd1e) $display("ERROR! at (14,16)\n");
if(PE_pixels_15_16!==16'h00e0) $display("ERROR! at (15,16)\n");
if(PE_pixels_16_16!==16'hf8cb) $display("ERROR! at (16,16)\n");
if(PE_pixels_17_16!==16'h00e1) $display("ERROR! at (17,16)\n");
if(PE_pixels_18_16!==16'h0064) $display("ERROR! at (18,16)\n");
if(PE_pixels_19_16!==16'h037a) $display("ERROR! at (19,16)\n");
if(PE_pixels_20_16!==16'hf7db) $display("ERROR! at (20,16)\n");
if(PE_pixels_21_16!==16'h0203) $display("ERROR! at (21,16)\n");
if(PE_pixels_22_16!==16'hfeb3) $display("ERROR! at (22,16)\n");
if(PE_pixels_23_16!==16'hff51) $display("ERROR! at (23,16)\n");
if(PE_pixels_24_16!==16'hfc71) $display("ERROR! at (24,16)\n");
if(PE_pixels_25_16!==16'hfe88) $display("ERROR! at (25,16)\n");
if(PE_pixels_26_16!==16'hfe53) $display("ERROR! at (26,16)\n");
if(PE_pixels_27_16!==16'h02d0) $display("ERROR! at (27,16)\n");
if(PE_pixels_28_16!==16'hfc9e) $display("ERROR! at (28,16)\n");
if(PE_pixels_29_16!==16'hfb77) $display("ERROR! at (29,16)\n");
if(PE_pixels_30_16!==16'h001f) $display("ERROR! at (30,16)\n");
if(PE_pixels_31_16!==16'h0066) $display("ERROR! at (31,16)\n");
if(PE_pixels_0_17!==16'h017c) $display("ERROR! at (0,17)\n");
if(PE_pixels_1_17!==16'hffb3) $display("ERROR! at (1,17)\n");
if(PE_pixels_2_17!==16'h008f) $display("ERROR! at (2,17)\n");
if(PE_pixels_3_17!==16'hfa1f) $display("ERROR! at (3,17)\n");
if(PE_pixels_4_17!==16'h0083) $display("ERROR! at (4,17)\n");
if(PE_pixels_5_17!==16'hffe2) $display("ERROR! at (5,17)\n");
if(PE_pixels_6_17!==16'h0504) $display("ERROR! at (6,17)\n");
if(PE_pixels_7_17!==16'hff3d) $display("ERROR! at (7,17)\n");
if(PE_pixels_8_17!==16'hfd82) $display("ERROR! at (8,17)\n");
if(PE_pixels_9_17!==16'h0083) $display("ERROR! at (9,17)\n");
if(PE_pixels_10_17!==16'hfe81) $display("ERROR! at (10,17)\n");
if(PE_pixels_11_17!==16'h02e3) $display("ERROR! at (11,17)\n");
if(PE_pixels_12_17!==16'h010f) $display("ERROR! at (12,17)\n");
if(PE_pixels_13_17!==16'h041b) $display("ERROR! at (13,17)\n");
if(PE_pixels_14_17!==16'h0203) $display("ERROR! at (14,17)\n");
if(PE_pixels_15_17!==16'hfd92) $display("ERROR! at (15,17)\n");
if(PE_pixels_16_17!==16'h007a) $display("ERROR! at (16,17)\n");
if(PE_pixels_17_17!==16'h0120) $display("ERROR! at (17,17)\n");
if(PE_pixels_18_17!==16'hfb0f) $display("ERROR! at (18,17)\n");
if(PE_pixels_19_17!==16'h013c) $display("ERROR! at (19,17)\n");
if(PE_pixels_20_17!==16'hfecc) $display("ERROR! at (20,17)\n");
if(PE_pixels_21_17!==16'hfd90) $display("ERROR! at (21,17)\n");
if(PE_pixels_22_17!==16'hff5f) $display("ERROR! at (22,17)\n");
if(PE_pixels_23_17!==16'h03d3) $display("ERROR! at (23,17)\n");
if(PE_pixels_24_17!==16'hfde9) $display("ERROR! at (24,17)\n");
if(PE_pixels_25_17!==16'h008e) $display("ERROR! at (25,17)\n");
if(PE_pixels_26_17!==16'hf92b) $display("ERROR! at (26,17)\n");
if(PE_pixels_27_17!==16'h025e) $display("ERROR! at (27,17)\n");
if(PE_pixels_28_17!==16'hf952) $display("ERROR! at (28,17)\n");
if(PE_pixels_29_17!==16'h046d) $display("ERROR! at (29,17)\n");
if(PE_pixels_30_17!==16'h012a) $display("ERROR! at (30,17)\n");
if(PE_pixels_31_17!==16'hff6d) $display("ERROR! at (31,17)\n");
if(PE_pixels_0_18!==16'h0036) $display("ERROR! at (0,18)\n");
if(PE_pixels_1_18!==16'h004e) $display("ERROR! at (1,18)\n");
if(PE_pixels_2_18!==16'hff97) $display("ERROR! at (2,18)\n");
if(PE_pixels_3_18!==16'hfe26) $display("ERROR! at (3,18)\n");
if(PE_pixels_4_18!==16'hfe8f) $display("ERROR! at (4,18)\n");
if(PE_pixels_5_18!==16'h018c) $display("ERROR! at (5,18)\n");
if(PE_pixels_6_18!==16'h05c6) $display("ERROR! at (6,18)\n");
if(PE_pixels_7_18!==16'hfd97) $display("ERROR! at (7,18)\n");
if(PE_pixels_8_18!==16'hff25) $display("ERROR! at (8,18)\n");
if(PE_pixels_9_18!==16'hfaef) $display("ERROR! at (9,18)\n");
if(PE_pixels_10_18!==16'hfdf7) $display("ERROR! at (10,18)\n");
if(PE_pixels_11_18!==16'hfda9) $display("ERROR! at (11,18)\n");
if(PE_pixels_12_18!==16'hfbc4) $display("ERROR! at (12,18)\n");
if(PE_pixels_13_18!==16'h07b2) $display("ERROR! at (13,18)\n");
if(PE_pixels_14_18!==16'hfe16) $display("ERROR! at (14,18)\n");
if(PE_pixels_15_18!==16'h06cd) $display("ERROR! at (15,18)\n");
if(PE_pixels_16_18!==16'hf592) $display("ERROR! at (16,18)\n");
if(PE_pixels_17_18!==16'hfd8b) $display("ERROR! at (17,18)\n");
if(PE_pixels_18_18!==16'hffcc) $display("ERROR! at (18,18)\n");
if(PE_pixels_19_18!==16'h0533) $display("ERROR! at (19,18)\n");
if(PE_pixels_20_18!==16'hfe4a) $display("ERROR! at (20,18)\n");
if(PE_pixels_21_18!==16'h017a) $display("ERROR! at (21,18)\n");
if(PE_pixels_22_18!==16'hfe31) $display("ERROR! at (22,18)\n");
if(PE_pixels_23_18!==16'h00e3) $display("ERROR! at (23,18)\n");
if(PE_pixels_24_18!==16'hffc9) $display("ERROR! at (24,18)\n");
if(PE_pixels_25_18!==16'h033e) $display("ERROR! at (25,18)\n");
if(PE_pixels_26_18!==16'h0236) $display("ERROR! at (26,18)\n");
if(PE_pixels_27_18!==16'h01d8) $display("ERROR! at (27,18)\n");
if(PE_pixels_28_18!==16'hfe6d) $display("ERROR! at (28,18)\n");
if(PE_pixels_29_18!==16'h01cf) $display("ERROR! at (29,18)\n");
if(PE_pixels_30_18!==16'hff07) $display("ERROR! at (30,18)\n");
if(PE_pixels_31_18!==16'hffc7) $display("ERROR! at (31,18)\n");
if(PE_pixels_0_19!==16'hff75) $display("ERROR! at (0,19)\n");
if(PE_pixels_1_19!==16'hffb8) $display("ERROR! at (1,19)\n");
if(PE_pixels_2_19!==16'hff0e) $display("ERROR! at (2,19)\n");
if(PE_pixels_3_19!==16'h0313) $display("ERROR! at (3,19)\n");
if(PE_pixels_4_19!==16'h009f) $display("ERROR! at (4,19)\n");
if(PE_pixels_5_19!==16'h01b2) $display("ERROR! at (5,19)\n");
if(PE_pixels_6_19!==16'hfbb7) $display("ERROR! at (6,19)\n");
if(PE_pixels_7_19!==16'hffb4) $display("ERROR! at (7,19)\n");
if(PE_pixels_8_19!==16'hfd77) $display("ERROR! at (8,19)\n");
if(PE_pixels_9_19!==16'hf952) $display("ERROR! at (9,19)\n");
if(PE_pixels_10_19!==16'hfee0) $display("ERROR! at (10,19)\n");
if(PE_pixels_11_19!==16'hfdc1) $display("ERROR! at (11,19)\n");
if(PE_pixels_12_19!==16'hfe59) $display("ERROR! at (12,19)\n");
if(PE_pixels_13_19!==16'h01cc) $display("ERROR! at (13,19)\n");
if(PE_pixels_14_19!==16'h024e) $display("ERROR! at (14,19)\n");
if(PE_pixels_15_19!==16'h036a) $display("ERROR! at (15,19)\n");
if(PE_pixels_16_19!==16'hfaa6) $display("ERROR! at (16,19)\n");
if(PE_pixels_17_19!==16'hfa1b) $display("ERROR! at (17,19)\n");
if(PE_pixels_18_19!==16'hfd8a) $display("ERROR! at (18,19)\n");
if(PE_pixels_19_19!==16'h0080) $display("ERROR! at (19,19)\n");
if(PE_pixels_20_19!==16'h085a) $display("ERROR! at (20,19)\n");
if(PE_pixels_21_19!==16'hff0d) $display("ERROR! at (21,19)\n");
if(PE_pixels_22_19!==16'hfbc0) $display("ERROR! at (22,19)\n");
if(PE_pixels_23_19!==16'h015e) $display("ERROR! at (23,19)\n");
if(PE_pixels_24_19!==16'h0030) $display("ERROR! at (24,19)\n");
if(PE_pixels_25_19!==16'h0382) $display("ERROR! at (25,19)\n");
if(PE_pixels_26_19!==16'hfd5b) $display("ERROR! at (26,19)\n");
if(PE_pixels_27_19!==16'hfc7b) $display("ERROR! at (27,19)\n");
if(PE_pixels_28_19!==16'hff64) $display("ERROR! at (28,19)\n");
if(PE_pixels_29_19!==16'h0030) $display("ERROR! at (29,19)\n");
if(PE_pixels_30_19!==16'h0018) $display("ERROR! at (30,19)\n");
if(PE_pixels_31_19!==16'hfd67) $display("ERROR! at (31,19)\n");
if(PE_pixels_0_20!==16'h00cb) $display("ERROR! at (0,20)\n");
if(PE_pixels_1_20!==16'h0016) $display("ERROR! at (1,20)\n");
if(PE_pixels_2_20!==16'hfdf7) $display("ERROR! at (2,20)\n");
if(PE_pixels_3_20!==16'h0079) $display("ERROR! at (3,20)\n");
if(PE_pixels_4_20!==16'hff8b) $display("ERROR! at (4,20)\n");
if(PE_pixels_5_20!==16'h0214) $display("ERROR! at (5,20)\n");
if(PE_pixels_6_20!==16'h067c) $display("ERROR! at (6,20)\n");
if(PE_pixels_7_20!==16'h0184) $display("ERROR! at (7,20)\n");
if(PE_pixels_8_20!==16'hfebc) $display("ERROR! at (8,20)\n");
if(PE_pixels_9_20!==16'hfe4f) $display("ERROR! at (9,20)\n");
if(PE_pixels_10_20!==16'hfc1e) $display("ERROR! at (10,20)\n");
if(PE_pixels_11_20!==16'h02ab) $display("ERROR! at (11,20)\n");
if(PE_pixels_12_20!==16'hf86a) $display("ERROR! at (12,20)\n");
if(PE_pixels_13_20!==16'hff75) $display("ERROR! at (13,20)\n");
if(PE_pixels_14_20!==16'hfc5a) $display("ERROR! at (14,20)\n");
if(PE_pixels_15_20!==16'h0796) $display("ERROR! at (15,20)\n");
if(PE_pixels_16_20!==16'h01b4) $display("ERROR! at (16,20)\n");
if(PE_pixels_17_20!==16'hfdd3) $display("ERROR! at (17,20)\n");
if(PE_pixels_18_20!==16'h029c) $display("ERROR! at (18,20)\n");
if(PE_pixels_19_20!==16'hfecc) $display("ERROR! at (19,20)\n");
if(PE_pixels_20_20!==16'h0188) $display("ERROR! at (20,20)\n");
if(PE_pixels_21_20!==16'hf79f) $display("ERROR! at (21,20)\n");
if(PE_pixels_22_20!==16'h0206) $display("ERROR! at (22,20)\n");
if(PE_pixels_23_20!==16'h0386) $display("ERROR! at (23,20)\n");
if(PE_pixels_24_20!==16'h0515) $display("ERROR! at (24,20)\n");
if(PE_pixels_25_20!==16'hfcf3) $display("ERROR! at (25,20)\n");
if(PE_pixels_26_20!==16'hfcc3) $display("ERROR! at (26,20)\n");
if(PE_pixels_27_20!==16'h00b3) $display("ERROR! at (27,20)\n");
if(PE_pixels_28_20!==16'hfd23) $display("ERROR! at (28,20)\n");
if(PE_pixels_29_20!==16'hfe68) $display("ERROR! at (29,20)\n");
if(PE_pixels_30_20!==16'hffe3) $display("ERROR! at (30,20)\n");
if(PE_pixels_31_20!==16'hfeaa) $display("ERROR! at (31,20)\n");
if(PE_pixels_0_21!==16'h0048) $display("ERROR! at (0,21)\n");
if(PE_pixels_1_21!==16'h00c8) $display("ERROR! at (1,21)\n");
if(PE_pixels_2_21!==16'hff3d) $display("ERROR! at (2,21)\n");
if(PE_pixels_3_21!==16'hfd89) $display("ERROR! at (3,21)\n");
if(PE_pixels_4_21!==16'hfd0d) $display("ERROR! at (4,21)\n");
if(PE_pixels_5_21!==16'h00cc) $display("ERROR! at (5,21)\n");
if(PE_pixels_6_21!==16'h01a6) $display("ERROR! at (6,21)\n");
if(PE_pixels_7_21!==16'h05a2) $display("ERROR! at (7,21)\n");
if(PE_pixels_8_21!==16'h02a2) $display("ERROR! at (8,21)\n");
if(PE_pixels_9_21!==16'h0101) $display("ERROR! at (9,21)\n");
if(PE_pixels_10_21!==16'hfaf4) $display("ERROR! at (10,21)\n");
if(PE_pixels_11_21!==16'hfdc4) $display("ERROR! at (11,21)\n");
if(PE_pixels_12_21!==16'hfda6) $display("ERROR! at (12,21)\n");
if(PE_pixels_13_21!==16'h0220) $display("ERROR! at (13,21)\n");
if(PE_pixels_14_21!==16'h01be) $display("ERROR! at (14,21)\n");
if(PE_pixels_15_21!==16'h033e) $display("ERROR! at (15,21)\n");
if(PE_pixels_16_21!==16'hff69) $display("ERROR! at (16,21)\n");
if(PE_pixels_17_21!==16'hfec0) $display("ERROR! at (17,21)\n");
if(PE_pixels_18_21!==16'hf59a) $display("ERROR! at (18,21)\n");
if(PE_pixels_19_21!==16'hfe90) $display("ERROR! at (19,21)\n");
if(PE_pixels_20_21!==16'hfcd7) $display("ERROR! at (20,21)\n");
if(PE_pixels_21_21!==16'hfdfe) $display("ERROR! at (21,21)\n");
if(PE_pixels_22_21!==16'hff39) $display("ERROR! at (22,21)\n");
if(PE_pixels_23_21!==16'h0239) $display("ERROR! at (23,21)\n");
if(PE_pixels_24_21!==16'hfe44) $display("ERROR! at (24,21)\n");
if(PE_pixels_25_21!==16'h01a5) $display("ERROR! at (25,21)\n");
if(PE_pixels_26_21!==16'h0268) $display("ERROR! at (26,21)\n");
if(PE_pixels_27_21!==16'hfb59) $display("ERROR! at (27,21)\n");
if(PE_pixels_28_21!==16'hfea1) $display("ERROR! at (28,21)\n");
if(PE_pixels_29_21!==16'hff00) $display("ERROR! at (29,21)\n");
if(PE_pixels_30_21!==16'h0312) $display("ERROR! at (30,21)\n");
if(PE_pixels_31_21!==16'hfea1) $display("ERROR! at (31,21)\n");
if(PE_pixels_0_22!==16'hff24) $display("ERROR! at (0,22)\n");
if(PE_pixels_1_22!==16'h0012) $display("ERROR! at (1,22)\n");
if(PE_pixels_2_22!==16'h01a7) $display("ERROR! at (2,22)\n");
if(PE_pixels_3_22!==16'h01bc) $display("ERROR! at (3,22)\n");
if(PE_pixels_4_22!==16'hfe68) $display("ERROR! at (4,22)\n");
if(PE_pixels_5_22!==16'hfbf0) $display("ERROR! at (5,22)\n");
if(PE_pixels_6_22!==16'hff80) $display("ERROR! at (6,22)\n");
if(PE_pixels_7_22!==16'h0222) $display("ERROR! at (7,22)\n");
if(PE_pixels_8_22!==16'h01a1) $display("ERROR! at (8,22)\n");
if(PE_pixels_9_22!==16'h00f2) $display("ERROR! at (9,22)\n");
if(PE_pixels_10_22!==16'hfbd4) $display("ERROR! at (10,22)\n");
if(PE_pixels_11_22!==16'hfeac) $display("ERROR! at (11,22)\n");
if(PE_pixels_12_22!==16'h00b7) $display("ERROR! at (12,22)\n");
if(PE_pixels_13_22!==16'h000b) $display("ERROR! at (13,22)\n");
if(PE_pixels_14_22!==16'h01c7) $display("ERROR! at (14,22)\n");
if(PE_pixels_15_22!==16'h00e8) $display("ERROR! at (15,22)\n");
if(PE_pixels_16_22!==16'h0554) $display("ERROR! at (16,22)\n");
if(PE_pixels_17_22!==16'hfced) $display("ERROR! at (17,22)\n");
if(PE_pixels_18_22!==16'hfdb1) $display("ERROR! at (18,22)\n");
if(PE_pixels_19_22!==16'hfe96) $display("ERROR! at (19,22)\n");
if(PE_pixels_20_22!==16'hfdea) $display("ERROR! at (20,22)\n");
if(PE_pixels_21_22!==16'hfcb9) $display("ERROR! at (21,22)\n");
if(PE_pixels_22_22!==16'hfb34) $display("ERROR! at (22,22)\n");
if(PE_pixels_23_22!==16'hfb0e) $display("ERROR! at (23,22)\n");
if(PE_pixels_24_22!==16'h00ff) $display("ERROR! at (24,22)\n");
if(PE_pixels_25_22!==16'h0016) $display("ERROR! at (25,22)\n");
if(PE_pixels_26_22!==16'hffc7) $display("ERROR! at (26,22)\n");
if(PE_pixels_27_22!==16'h0678) $display("ERROR! at (27,22)\n");
if(PE_pixels_28_22!==16'h00e5) $display("ERROR! at (28,22)\n");
if(PE_pixels_29_22!==16'hfec9) $display("ERROR! at (29,22)\n");
if(PE_pixels_30_22!==16'hffdd) $display("ERROR! at (30,22)\n");
if(PE_pixels_31_22!==16'hfcf3) $display("ERROR! at (31,22)\n");
if(PE_pixels_0_23!==16'hff7c) $display("ERROR! at (0,23)\n");
if(PE_pixels_1_23!==16'h011d) $display("ERROR! at (1,23)\n");
if(PE_pixels_2_23!==16'h0230) $display("ERROR! at (2,23)\n");
if(PE_pixels_3_23!==16'h0270) $display("ERROR! at (3,23)\n");
if(PE_pixels_4_23!==16'hfeb4) $display("ERROR! at (4,23)\n");
if(PE_pixels_5_23!==16'hfb82) $display("ERROR! at (5,23)\n");
if(PE_pixels_6_23!==16'h018f) $display("ERROR! at (6,23)\n");
if(PE_pixels_7_23!==16'hfd5e) $display("ERROR! at (7,23)\n");
if(PE_pixels_8_23!==16'h0023) $display("ERROR! at (8,23)\n");
if(PE_pixels_9_23!==16'h0114) $display("ERROR! at (9,23)\n");
if(PE_pixels_10_23!==16'hfd05) $display("ERROR! at (10,23)\n");
if(PE_pixels_11_23!==16'hfbbf) $display("ERROR! at (11,23)\n");
if(PE_pixels_12_23!==16'h001c) $display("ERROR! at (12,23)\n");
if(PE_pixels_13_23!==16'hff46) $display("ERROR! at (13,23)\n");
if(PE_pixels_14_23!==16'hfe74) $display("ERROR! at (14,23)\n");
if(PE_pixels_15_23!==16'hfd56) $display("ERROR! at (15,23)\n");
if(PE_pixels_16_23!==16'h00e4) $display("ERROR! at (16,23)\n");
if(PE_pixels_17_23!==16'h0596) $display("ERROR! at (17,23)\n");
if(PE_pixels_18_23!==16'hfb74) $display("ERROR! at (18,23)\n");
if(PE_pixels_19_23!==16'h041d) $display("ERROR! at (19,23)\n");
if(PE_pixels_20_23!==16'h047f) $display("ERROR! at (20,23)\n");
if(PE_pixels_21_23!==16'hffa1) $display("ERROR! at (21,23)\n");
if(PE_pixels_22_23!==16'hf8a9) $display("ERROR! at (22,23)\n");
if(PE_pixels_23_23!==16'hf895) $display("ERROR! at (23,23)\n");
if(PE_pixels_24_23!==16'hfcb9) $display("ERROR! at (24,23)\n");
if(PE_pixels_25_23!==16'h0068) $display("ERROR! at (25,23)\n");
if(PE_pixels_26_23!==16'h08f3) $display("ERROR! at (26,23)\n");
if(PE_pixels_27_23!==16'hfef4) $display("ERROR! at (27,23)\n");
if(PE_pixels_28_23!==16'h00e3) $display("ERROR! at (28,23)\n");
if(PE_pixels_29_23!==16'h043a) $display("ERROR! at (29,23)\n");
if(PE_pixels_30_23!==16'hfd5d) $display("ERROR! at (30,23)\n");
if(PE_pixels_31_23!==16'hff28) $display("ERROR! at (31,23)\n");
if(PE_pixels_0_24!==16'hfe58) $display("ERROR! at (0,24)\n");
if(PE_pixels_1_24!==16'h00bb) $display("ERROR! at (1,24)\n");
if(PE_pixels_2_24!==16'h0171) $display("ERROR! at (2,24)\n");
if(PE_pixels_3_24!==16'h0165) $display("ERROR! at (3,24)\n");
if(PE_pixels_4_24!==16'h02b5) $display("ERROR! at (4,24)\n");
if(PE_pixels_5_24!==16'h0120) $display("ERROR! at (5,24)\n");
if(PE_pixels_6_24!==16'h01bd) $display("ERROR! at (6,24)\n");
if(PE_pixels_7_24!==16'h0045) $display("ERROR! at (7,24)\n");
if(PE_pixels_8_24!==16'h0180) $display("ERROR! at (8,24)\n");
if(PE_pixels_9_24!==16'hfc48) $display("ERROR! at (9,24)\n");
if(PE_pixels_10_24!==16'hfcf2) $display("ERROR! at (10,24)\n");
if(PE_pixels_11_24!==16'hfd4d) $display("ERROR! at (11,24)\n");
if(PE_pixels_12_24!==16'hfe32) $display("ERROR! at (12,24)\n");
if(PE_pixels_13_24!==16'h01c6) $display("ERROR! at (13,24)\n");
if(PE_pixels_14_24!==16'hff92) $display("ERROR! at (14,24)\n");
if(PE_pixels_15_24!==16'h0321) $display("ERROR! at (15,24)\n");
if(PE_pixels_16_24!==16'h0374) $display("ERROR! at (16,24)\n");
if(PE_pixels_17_24!==16'hff36) $display("ERROR! at (17,24)\n");
if(PE_pixels_18_24!==16'hfb65) $display("ERROR! at (18,24)\n");
if(PE_pixels_19_24!==16'hfd1a) $display("ERROR! at (19,24)\n");
if(PE_pixels_20_24!==16'h03fd) $display("ERROR! at (20,24)\n");
if(PE_pixels_21_24!==16'h061b) $display("ERROR! at (21,24)\n");
if(PE_pixels_22_24!==16'h0322) $display("ERROR! at (22,24)\n");
if(PE_pixels_23_24!==16'hf4a1) $display("ERROR! at (23,24)\n");
if(PE_pixels_24_24!==16'hfbe2) $display("ERROR! at (24,24)\n");
if(PE_pixels_25_24!==16'hfec9) $display("ERROR! at (25,24)\n");
if(PE_pixels_26_24!==16'hfe43) $display("ERROR! at (26,24)\n");
if(PE_pixels_27_24!==16'h010f) $display("ERROR! at (27,24)\n");
if(PE_pixels_28_24!==16'h040c) $display("ERROR! at (28,24)\n");
if(PE_pixels_29_24!==16'h00f2) $display("ERROR! at (29,24)\n");
if(PE_pixels_30_24!==16'h016e) $display("ERROR! at (30,24)\n");
if(PE_pixels_31_24!==16'hff04) $display("ERROR! at (31,24)\n");
if(PE_pixels_0_25!==16'hfdf8) $display("ERROR! at (0,25)\n");
if(PE_pixels_1_25!==16'hfffe) $display("ERROR! at (1,25)\n");
if(PE_pixels_2_25!==16'h0192) $display("ERROR! at (2,25)\n");
if(PE_pixels_3_25!==16'h0250) $display("ERROR! at (3,25)\n");
if(PE_pixels_4_25!==16'h06be) $display("ERROR! at (4,25)\n");
if(PE_pixels_5_25!==16'h00f4) $display("ERROR! at (5,25)\n");
if(PE_pixels_6_25!==16'h032e) $display("ERROR! at (6,25)\n");
if(PE_pixels_7_25!==16'h0061) $display("ERROR! at (7,25)\n");
if(PE_pixels_8_25!==16'h024f) $display("ERROR! at (8,25)\n");
if(PE_pixels_9_25!==16'h01e1) $display("ERROR! at (9,25)\n");
if(PE_pixels_10_25!==16'h0541) $display("ERROR! at (10,25)\n");
if(PE_pixels_11_25!==16'hfbe9) $display("ERROR! at (11,25)\n");
if(PE_pixels_12_25!==16'hfb15) $display("ERROR! at (12,25)\n");
if(PE_pixels_13_25!==16'hfdd0) $display("ERROR! at (13,25)\n");
if(PE_pixels_14_25!==16'h028a) $display("ERROR! at (14,25)\n");
if(PE_pixels_15_25!==16'h00bb) $display("ERROR! at (15,25)\n");
if(PE_pixels_16_25!==16'h015e) $display("ERROR! at (16,25)\n");
if(PE_pixels_17_25!==16'h0022) $display("ERROR! at (17,25)\n");
if(PE_pixels_18_25!==16'h001f) $display("ERROR! at (18,25)\n");
if(PE_pixels_19_25!==16'hfef4) $display("ERROR! at (19,25)\n");
if(PE_pixels_20_25!==16'hfc7f) $display("ERROR! at (20,25)\n");
if(PE_pixels_21_25!==16'h053f) $display("ERROR! at (21,25)\n");
if(PE_pixels_22_25!==16'hfd6c) $display("ERROR! at (22,25)\n");
if(PE_pixels_23_25!==16'h0159) $display("ERROR! at (23,25)\n");
if(PE_pixels_24_25!==16'hf757) $display("ERROR! at (24,25)\n");
if(PE_pixels_25_25!==16'h00ed) $display("ERROR! at (25,25)\n");
if(PE_pixels_26_25!==16'h01a9) $display("ERROR! at (26,25)\n");
if(PE_pixels_27_25!==16'hffec) $display("ERROR! at (27,25)\n");
if(PE_pixels_28_25!==16'hfc2e) $display("ERROR! at (28,25)\n");
if(PE_pixels_29_25!==16'h03ac) $display("ERROR! at (29,25)\n");
if(PE_pixels_30_25!==16'h0062) $display("ERROR! at (30,25)\n");
if(PE_pixels_31_25!==16'hff1c) $display("ERROR! at (31,25)\n");
if(PE_pixels_0_26!==16'hfe88) $display("ERROR! at (0,26)\n");
if(PE_pixels_1_26!==16'hff63) $display("ERROR! at (1,26)\n");
if(PE_pixels_2_26!==16'h01c1) $display("ERROR! at (2,26)\n");
if(PE_pixels_3_26!==16'hfe0a) $display("ERROR! at (3,26)\n");
if(PE_pixels_4_26!==16'h081c) $display("ERROR! at (4,26)\n");
if(PE_pixels_5_26!==16'h01b0) $display("ERROR! at (5,26)\n");
if(PE_pixels_6_26!==16'h0128) $display("ERROR! at (6,26)\n");
if(PE_pixels_7_26!==16'hfe6a) $display("ERROR! at (7,26)\n");
if(PE_pixels_8_26!==16'h0186) $display("ERROR! at (8,26)\n");
if(PE_pixels_9_26!==16'h0235) $display("ERROR! at (9,26)\n");
if(PE_pixels_10_26!==16'h0480) $display("ERROR! at (10,26)\n");
if(PE_pixels_11_26!==16'hfc15) $display("ERROR! at (11,26)\n");
if(PE_pixels_12_26!==16'hff9f) $display("ERROR! at (12,26)\n");
if(PE_pixels_13_26!==16'hff3f) $display("ERROR! at (13,26)\n");
if(PE_pixels_14_26!==16'hfea1) $display("ERROR! at (14,26)\n");
if(PE_pixels_15_26!==16'hfef0) $display("ERROR! at (15,26)\n");
if(PE_pixels_16_26!==16'hfc05) $display("ERROR! at (16,26)\n");
if(PE_pixels_17_26!==16'h0108) $display("ERROR! at (17,26)\n");
if(PE_pixels_18_26!==16'hfd5d) $display("ERROR! at (18,26)\n");
if(PE_pixels_19_26!==16'hfc10) $display("ERROR! at (19,26)\n");
if(PE_pixels_20_26!==16'hfcf6) $display("ERROR! at (20,26)\n");
if(PE_pixels_21_26!==16'h00e3) $display("ERROR! at (21,26)\n");
if(PE_pixels_22_26!==16'h0445) $display("ERROR! at (22,26)\n");
if(PE_pixels_23_26!==16'h0a8b) $display("ERROR! at (23,26)\n");
if(PE_pixels_24_26!==16'hfa01) $display("ERROR! at (24,26)\n");
if(PE_pixels_25_26!==16'hffb2) $display("ERROR! at (25,26)\n");
if(PE_pixels_26_26!==16'hfb2c) $display("ERROR! at (26,26)\n");
if(PE_pixels_27_26!==16'hff53) $display("ERROR! at (27,26)\n");
if(PE_pixels_28_26!==16'hffd6) $display("ERROR! at (28,26)\n");
if(PE_pixels_29_26!==16'h01c9) $display("ERROR! at (29,26)\n");
if(PE_pixels_30_26!==16'hfe45) $display("ERROR! at (30,26)\n");
if(PE_pixels_31_26!==16'hffb0) $display("ERROR! at (31,26)\n");
if(PE_pixels_0_27!==16'h0062) $display("ERROR! at (0,27)\n");
if(PE_pixels_1_27!==16'hfc78) $display("ERROR! at (1,27)\n");
if(PE_pixels_2_27!==16'hfec2) $display("ERROR! at (2,27)\n");
if(PE_pixels_3_27!==16'h0133) $display("ERROR! at (3,27)\n");
if(PE_pixels_4_27!==16'h0845) $display("ERROR! at (4,27)\n");
if(PE_pixels_5_27!==16'hff81) $display("ERROR! at (5,27)\n");
if(PE_pixels_6_27!==16'hfa4b) $display("ERROR! at (6,27)\n");
if(PE_pixels_7_27!==16'h01e2) $display("ERROR! at (7,27)\n");
if(PE_pixels_8_27!==16'hfa84) $display("ERROR! at (8,27)\n");
if(PE_pixels_9_27!==16'h0220) $display("ERROR! at (9,27)\n");
if(PE_pixels_10_27!==16'h0161) $display("ERROR! at (10,27)\n");
if(PE_pixels_11_27!==16'h0261) $display("ERROR! at (11,27)\n");
if(PE_pixels_12_27!==16'hfd7c) $display("ERROR! at (12,27)\n");
if(PE_pixels_13_27!==16'h024d) $display("ERROR! at (13,27)\n");
if(PE_pixels_14_27!==16'hfdca) $display("ERROR! at (14,27)\n");
if(PE_pixels_15_27!==16'h0116) $display("ERROR! at (15,27)\n");
if(PE_pixels_16_27!==16'hfb3f) $display("ERROR! at (16,27)\n");
if(PE_pixels_17_27!==16'hfa48) $display("ERROR! at (17,27)\n");
if(PE_pixels_18_27!==16'hfcfd) $display("ERROR! at (18,27)\n");
if(PE_pixels_19_27!==16'hfffc) $display("ERROR! at (19,27)\n");
if(PE_pixels_20_27!==16'hf8fe) $display("ERROR! at (20,27)\n");
if(PE_pixels_21_27!==16'hff03) $display("ERROR! at (21,27)\n");
if(PE_pixels_22_27!==16'h03fb) $display("ERROR! at (22,27)\n");
if(PE_pixels_23_27!==16'h0652) $display("ERROR! at (23,27)\n");
if(PE_pixels_24_27!==16'hff12) $display("ERROR! at (24,27)\n");
if(PE_pixels_25_27!==16'hfda4) $display("ERROR! at (25,27)\n");
if(PE_pixels_26_27!==16'h01dc) $display("ERROR! at (26,27)\n");
if(PE_pixels_27_27!==16'hfd26) $display("ERROR! at (27,27)\n");
if(PE_pixels_28_27!==16'h01a8) $display("ERROR! at (28,27)\n");
if(PE_pixels_29_27!==16'h01d7) $display("ERROR! at (29,27)\n");
if(PE_pixels_30_27!==16'hff09) $display("ERROR! at (30,27)\n");
if(PE_pixels_31_27!==16'h02d8) $display("ERROR! at (31,27)\n");
if(PE_pixels_0_28!==16'h0261) $display("ERROR! at (0,28)\n");
if(PE_pixels_1_28!==16'hfec9) $display("ERROR! at (1,28)\n");
if(PE_pixels_2_28!==16'h010e) $display("ERROR! at (2,28)\n");
if(PE_pixels_3_28!==16'hfb78) $display("ERROR! at (3,28)\n");
if(PE_pixels_4_28!==16'h02c2) $display("ERROR! at (4,28)\n");
if(PE_pixels_5_28!==16'h01b0) $display("ERROR! at (5,28)\n");
if(PE_pixels_6_28!==16'hfb8c) $display("ERROR! at (6,28)\n");
if(PE_pixels_7_28!==16'h01f7) $display("ERROR! at (7,28)\n");
if(PE_pixels_8_28!==16'hfac7) $display("ERROR! at (8,28)\n");
if(PE_pixels_9_28!==16'h0132) $display("ERROR! at (9,28)\n");
if(PE_pixels_10_28!==16'h000a) $display("ERROR! at (10,28)\n");
if(PE_pixels_11_28!==16'h02ce) $display("ERROR! at (11,28)\n");
if(PE_pixels_12_28!==16'hfbd8) $display("ERROR! at (12,28)\n");
if(PE_pixels_13_28!==16'h0089) $display("ERROR! at (13,28)\n");
if(PE_pixels_14_28!==16'h0240) $display("ERROR! at (14,28)\n");
if(PE_pixels_15_28!==16'h0202) $display("ERROR! at (15,28)\n");
if(PE_pixels_16_28!==16'hfd74) $display("ERROR! at (16,28)\n");
if(PE_pixels_17_28!==16'hfd7e) $display("ERROR! at (17,28)\n");
if(PE_pixels_18_28!==16'hfcf9) $display("ERROR! at (18,28)\n");
if(PE_pixels_19_28!==16'h00ee) $display("ERROR! at (19,28)\n");
if(PE_pixels_20_28!==16'h04f9) $display("ERROR! at (20,28)\n");
if(PE_pixels_21_28!==16'hfe39) $display("ERROR! at (21,28)\n");
if(PE_pixels_22_28!==16'hfc9b) $display("ERROR! at (22,28)\n");
if(PE_pixels_23_28!==16'hff69) $display("ERROR! at (23,28)\n");
if(PE_pixels_24_28!==16'h02b1) $display("ERROR! at (24,28)\n");
if(PE_pixels_25_28!==16'h0040) $display("ERROR! at (25,28)\n");
if(PE_pixels_26_28!==16'hfaa7) $display("ERROR! at (26,28)\n");
if(PE_pixels_27_28!==16'h02f6) $display("ERROR! at (27,28)\n");
if(PE_pixels_28_28!==16'hfb14) $display("ERROR! at (28,28)\n");
if(PE_pixels_29_28!==16'h044d) $display("ERROR! at (29,28)\n");
if(PE_pixels_30_28!==16'h0414) $display("ERROR! at (30,28)\n");
if(PE_pixels_31_28!==16'h0073) $display("ERROR! at (31,28)\n");
if(PE_pixels_0_29!==16'hffdb) $display("ERROR! at (0,29)\n");
if(PE_pixels_1_29!==16'hfe5d) $display("ERROR! at (1,29)\n");
if(PE_pixels_2_29!==16'hfd71) $display("ERROR! at (2,29)\n");
if(PE_pixels_3_29!==16'hffd1) $display("ERROR! at (3,29)\n");
if(PE_pixels_4_29!==16'h0077) $display("ERROR! at (4,29)\n");
if(PE_pixels_5_29!==16'h005d) $display("ERROR! at (5,29)\n");
if(PE_pixels_6_29!==16'hfedd) $display("ERROR! at (6,29)\n");
if(PE_pixels_7_29!==16'h09c5) $display("ERROR! at (7,29)\n");
if(PE_pixels_8_29!==16'hfa8a) $display("ERROR! at (8,29)\n");
if(PE_pixels_9_29!==16'h00b2) $display("ERROR! at (9,29)\n");
if(PE_pixels_10_29!==16'hfc5c) $display("ERROR! at (10,29)\n");
if(PE_pixels_11_29!==16'h0252) $display("ERROR! at (11,29)\n");
if(PE_pixels_12_29!==16'h008e) $display("ERROR! at (12,29)\n");
if(PE_pixels_13_29!==16'hfed6) $display("ERROR! at (13,29)\n");
if(PE_pixels_14_29!==16'hf9a3) $display("ERROR! at (14,29)\n");
if(PE_pixels_15_29!==16'h00a6) $display("ERROR! at (15,29)\n");
if(PE_pixels_16_29!==16'h03f4) $display("ERROR! at (16,29)\n");
if(PE_pixels_17_29!==16'h02c5) $display("ERROR! at (17,29)\n");
if(PE_pixels_18_29!==16'hfdef) $display("ERROR! at (18,29)\n");
if(PE_pixels_19_29!==16'h01eb) $display("ERROR! at (19,29)\n");
if(PE_pixels_20_29!==16'h0182) $display("ERROR! at (20,29)\n");
if(PE_pixels_21_29!==16'hfd59) $display("ERROR! at (21,29)\n");
if(PE_pixels_22_29!==16'h01b8) $display("ERROR! at (22,29)\n");
if(PE_pixels_23_29!==16'hfb4c) $display("ERROR! at (23,29)\n");
if(PE_pixels_24_29!==16'hffd0) $display("ERROR! at (24,29)\n");
if(PE_pixels_25_29!==16'hfef5) $display("ERROR! at (25,29)\n");
if(PE_pixels_26_29!==16'h04c0) $display("ERROR! at (26,29)\n");
if(PE_pixels_27_29!==16'hfec7) $display("ERROR! at (27,29)\n");
if(PE_pixels_28_29!==16'hfeb1) $display("ERROR! at (28,29)\n");
if(PE_pixels_29_29!==16'h03e5) $display("ERROR! at (29,29)\n");
if(PE_pixels_30_29!==16'hfd19) $display("ERROR! at (30,29)\n");
if(PE_pixels_31_29!==16'h0126) $display("ERROR! at (31,29)\n");
if(PE_pixels_0_30!==16'h0000) $display("ERROR! at (0,30)\n");
if(PE_pixels_1_30!==16'h0088) $display("ERROR! at (1,30)\n");
if(PE_pixels_2_30!==16'hff67) $display("ERROR! at (2,30)\n");
if(PE_pixels_3_30!==16'h0050) $display("ERROR! at (3,30)\n");
if(PE_pixels_4_30!==16'hfe8a) $display("ERROR! at (4,30)\n");
if(PE_pixels_5_30!==16'h036a) $display("ERROR! at (5,30)\n");
if(PE_pixels_6_30!==16'hffd4) $display("ERROR! at (6,30)\n");
if(PE_pixels_7_30!==16'hff8d) $display("ERROR! at (7,30)\n");
if(PE_pixels_8_30!==16'hfc12) $display("ERROR! at (8,30)\n");
if(PE_pixels_9_30!==16'h029f) $display("ERROR! at (9,30)\n");
if(PE_pixels_10_30!==16'hfea3) $display("ERROR! at (10,30)\n");
if(PE_pixels_11_30!==16'hff44) $display("ERROR! at (11,30)\n");
if(PE_pixels_12_30!==16'h0151) $display("ERROR! at (12,30)\n");
if(PE_pixels_13_30!==16'hff09) $display("ERROR! at (13,30)\n");
if(PE_pixels_14_30!==16'h06c9) $display("ERROR! at (14,30)\n");
if(PE_pixels_15_30!==16'hfec9) $display("ERROR! at (15,30)\n");
if(PE_pixels_16_30!==16'h02d6) $display("ERROR! at (16,30)\n");
if(PE_pixels_17_30!==16'hfe16) $display("ERROR! at (17,30)\n");
if(PE_pixels_18_30!==16'hfd11) $display("ERROR! at (18,30)\n");
if(PE_pixels_19_30!==16'h0069) $display("ERROR! at (19,30)\n");
if(PE_pixels_20_30!==16'hff6e) $display("ERROR! at (20,30)\n");
if(PE_pixels_21_30!==16'hfdd1) $display("ERROR! at (21,30)\n");
if(PE_pixels_22_30!==16'hfe25) $display("ERROR! at (22,30)\n");
if(PE_pixels_23_30!==16'h020b) $display("ERROR! at (23,30)\n");
if(PE_pixels_24_30!==16'h0343) $display("ERROR! at (24,30)\n");
if(PE_pixels_25_30!==16'h00c1) $display("ERROR! at (25,30)\n");
if(PE_pixels_26_30!==16'hfd21) $display("ERROR! at (26,30)\n");
if(PE_pixels_27_30!==16'h0403) $display("ERROR! at (27,30)\n");
if(PE_pixels_28_30!==16'hfe9f) $display("ERROR! at (28,30)\n");
if(PE_pixels_29_30!==16'hf966) $display("ERROR! at (29,30)\n");
if(PE_pixels_30_30!==16'h0391) $display("ERROR! at (30,30)\n");
if(PE_pixels_31_30!==16'h00e9) $display("ERROR! at (31,30)\n");
if(PE_pixels_0_31!==16'h0000) $display("ERROR! at (0,31)\n");
if(PE_pixels_1_31!==16'hfff8) $display("ERROR! at (1,31)\n");
if(PE_pixels_2_31!==16'hffb9) $display("ERROR! at (2,31)\n");
if(PE_pixels_3_31!==16'hffe2) $display("ERROR! at (3,31)\n");
if(PE_pixels_4_31!==16'h006f) $display("ERROR! at (4,31)\n");
if(PE_pixels_5_31!==16'h00b3) $display("ERROR! at (5,31)\n");
if(PE_pixels_6_31!==16'hff64) $display("ERROR! at (6,31)\n");
if(PE_pixels_7_31!==16'h0096) $display("ERROR! at (7,31)\n");
if(PE_pixels_8_31!==16'h00e1) $display("ERROR! at (8,31)\n");
if(PE_pixels_9_31!==16'h002d) $display("ERROR! at (9,31)\n");
if(PE_pixels_10_31!==16'hfee3) $display("ERROR! at (10,31)\n");
if(PE_pixels_11_31!==16'h001c) $display("ERROR! at (11,31)\n");
if(PE_pixels_12_31!==16'h0104) $display("ERROR! at (12,31)\n");
if(PE_pixels_13_31!==16'h00dc) $display("ERROR! at (13,31)\n");
if(PE_pixels_14_31!==16'hff28) $display("ERROR! at (14,31)\n");
if(PE_pixels_15_31!==16'hfdab) $display("ERROR! at (15,31)\n");
if(PE_pixels_16_31!==16'h014a) $display("ERROR! at (16,31)\n");
if(PE_pixels_17_31!==16'hffb5) $display("ERROR! at (17,31)\n");
if(PE_pixels_18_31!==16'hfff1) $display("ERROR! at (18,31)\n");
if(PE_pixels_19_31!==16'h005f) $display("ERROR! at (19,31)\n");
if(PE_pixels_20_31!==16'h0007) $display("ERROR! at (20,31)\n");
if(PE_pixels_21_31!==16'h0057) $display("ERROR! at (21,31)\n");
if(PE_pixels_22_31!==16'h0113) $display("ERROR! at (22,31)\n");
if(PE_pixels_23_31!==16'h00f8) $display("ERROR! at (23,31)\n");
if(PE_pixels_24_31!==16'hfead) $display("ERROR! at (24,31)\n");
if(PE_pixels_25_31!==16'hfdff) $display("ERROR! at (25,31)\n");
if(PE_pixels_26_31!==16'h00e4) $display("ERROR! at (26,31)\n");
if(PE_pixels_27_31!==16'h0116) $display("ERROR! at (27,31)\n");
if(PE_pixels_28_31!==16'hfca2) $display("ERROR! at (28,31)\n");
if(PE_pixels_29_31!==16'h0006) $display("ERROR! at (29,31)\n");
if(PE_pixels_30_31!==16'h0288) $display("ERROR! at (30,31)\n");
if(PE_pixels_31_31!==16'hff7b) $display("ERROR! at (31,31)\n");






    $finish;
    
end
reg test_valid;
always@(posedge clk)begin
    if(rst)begin
        test_valid<= 'd0;
    end
    else begin
        test_valid = CSR_valid;
        if(PE_out_valid)begin
            
            PE_result[ (($signed(PE_col_answer_1_1)+4)+($signed(PE_row_answer_1_1)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_1_1)+4)+($signed(PE_row_answer_1_1)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_1_1);
            PE_result[ (($signed(PE_col_answer_1_2)+4)+($signed(PE_row_answer_1_2)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_1_2)+4)+($signed(PE_row_answer_1_2)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_1_2);
            PE_result[ (($signed(PE_col_answer_1_3)+4)+($signed(PE_row_answer_1_3)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_1_3)+4)+($signed(PE_row_answer_1_3)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_1_3);
            PE_result[ (($signed(PE_col_answer_1_4)+4)+($signed(PE_row_answer_1_4)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_1_4)+4)+($signed(PE_row_answer_1_4)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_1_4);

            PE_result[ (($signed(PE_col_answer_2_1)+4)+($signed(PE_row_answer_2_1)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_2_1)+4)+($signed(PE_row_answer_2_1)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_2_1);
            PE_result[ (($signed(PE_col_answer_2_2)+4)+($signed(PE_row_answer_2_2)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_2_2)+4)+($signed(PE_row_answer_2_2)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_2_2);
            PE_result[ (($signed(PE_col_answer_2_3)+4)+($signed(PE_row_answer_2_3)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_2_3)+4)+($signed(PE_row_answer_2_3)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_2_3);
            PE_result[ (($signed(PE_col_answer_2_4)+4)+($signed(PE_row_answer_2_4)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_2_4)+4)+($signed(PE_row_answer_2_4)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_2_4);

            PE_result[ (($signed(PE_col_answer_3_1)+4)+($signed(PE_row_answer_3_1)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_3_1)+4)+($signed(PE_row_answer_3_1)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_3_1);
            PE_result[ (($signed(PE_col_answer_3_2)+4)+($signed(PE_row_answer_3_2)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_3_2)+4)+($signed(PE_row_answer_3_2)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_3_2);
            PE_result[ (($signed(PE_col_answer_3_3)+4)+($signed(PE_row_answer_3_3)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_3_3)+4)+($signed(PE_row_answer_3_3)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_3_3);
            PE_result[ (($signed(PE_col_answer_3_4)+4)+($signed(PE_row_answer_3_4)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_3_4)+4)+($signed(PE_row_answer_3_4)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_3_4);

            PE_result[ (($signed(PE_col_answer_4_1)+4)+($signed(PE_row_answer_4_1)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_4_1)+4)+($signed(PE_row_answer_4_1)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_4_1);
            PE_result[ (($signed(PE_col_answer_4_2)+4)+($signed(PE_row_answer_4_2)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_4_2)+4)+($signed(PE_row_answer_4_2)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_4_2);
            PE_result[ (($signed(PE_col_answer_4_3)+4)+($signed(PE_row_answer_4_3)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_4_3)+4)+($signed(PE_row_answer_4_3)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_4_3);
            PE_result[ (($signed(PE_col_answer_4_4)+4)+($signed(PE_row_answer_4_4)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(PE_result[ (($signed(PE_col_answer_4_4)+4)+($signed(PE_row_answer_4_4)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(PE_answer_4_4);

        end 
    end

    //PE_result[11*(data_out_rows[col_length-1:0]+4)+(data_out_cols[col_length-1:0]+4)+1 -:word_length] <= data_out[word_length-1:0] + PE_result[11*(data_out_rows[col_length-1:0]+4)+(data_out_cols[col_length-1:0]+4)+1 -:word_length];
end



always #5 clk = ~clk;
CSR#
(
    .col_length(col_length), 
    .word_length(word_length), 
    .double_word_length(double_word_length), 
    .kernel_size(kernel_size), 
    .image_size(image_size)
)u1
(
    .clk(clk), 
    .rst(rst), 
    .in_valid(in_valid),
    .data_in(data_in),
    .data_out(CSR_data_out),
    .data_out_cols(CSR_data_out_cols),
    .data_out_rows(CSR_data_out_rows),
    .valid_num_out(valid_num_out),
    .out_valid(CSR_valid)
);

PE#
(
    .col_length(col_length), 
    .word_length(word_length), 
    .double_word_length(double_word_length), 
    .kernel_size(kernel_size), 
    .image_size(image_size)
)u2
(
    .clk(clk), 
    .rst(rst), 
    .in_valid(CSR_valid),
    .in_channel(in_channel),
    .feature_valid_num(valid_num_out),
    .feature_value(CSR_data_out),
    .feature_cols(CSR_data_out_cols),
    .feature_rows(CSR_data_out_rows),
    .weight_valid_num(weight_valid_num),
    .weight_value(pe_input_weight_value),
    .weight_cols(pe_input_weight_cols),
    .weight_rows(pe_input_weight_rows),
    .data_out(PE_data_out),
    .data_out_cols(PE_data_out_cols),
    .data_out_rows(PE_data_out_rows),
    .out_valid(PE_out_valid),
    .out_channel(out_channel)
);



endmodule