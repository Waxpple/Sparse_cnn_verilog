`timescale 1ns/1ns
module CSR_tb();
parameter col_length = 8;
parameter word_length = 8;
parameter double_word_length = 16;
parameter kernel_size = 5;
parameter image_size = 36;

reg clk;
reg rst;
reg signed [word_length-1:0] data_in;
reg in_valid;
reg [10368-1 :0] pe_input_feature_value='h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_f0_dd_39_f3_f7_06_02_f7_02_f6_fc_15_f9_ff_15_08_fe_fb_f0_01_e5_09_00_f9_1d_fa_f6_ec_00_00_00_00_00_00_00_00_fd_f2_fb_f2_eb_f3_fa_f3_12_fc_f8_0b_03_fe_f1_f6_07_f7_eb_0a_17_f5_05_01_18_1f_f1_09_00_00_00_00_00_00_00_00_07_04_f3_0c_fa_f6_01_0d_07_e5_06_f8_0e_0b_f9_03_fc_e1_0b_f2_15_fa_0d_ee_08_f9_ed_ff_00_00_00_00_00_00_00_00_f8_fc_fa_f8_e8_07_f2_0f_00_da_08_fb_03_06_f2_f0_07_03_06_fb_e9_f5_13_06_fa_0d_05_0a_00_00_00_00_00_00_00_00_f1_0d_f6_03_fa_03_17_1c_06_e4_13_03_11_0c_f4_15_fb_0d_fd_07_02_0b_f5_0e_ea_e0_ee_04_00_00_00_00_00_00_00_00_f2_fb_01_01_e7_01_ea_07_0e_fc_08_1f_1a_04_fa_ef_02_00_d8_fa_eb_ee_0d_f1_f4_ff_01_fd_00_00_00_00_00_00_00_00_18_eb_f2_08_12_04_0b_fb_f7_0a_00_0b_05_f7_f2_0a_1a_e6_15_0e_29_12_f8_08_dd_f9_0f_10_00_00_00_00_00_00_00_00_05_df_02_07_f1_fe_01_0c_dc_fb_fb_fb_16_15_e8_f8_02_fe_0e_10_0d_fb_fa_02_fd_e5_03_09_00_00_00_00_00_00_00_00_f5_f9_fd_e5_05_0a_03_04_0c_0a_1d_0f_0e_1b_fb_26_f2_ec_08_08_f8_03_08_1b_fc_19_f7_f4_00_00_00_00_00_00_00_00_13_00_fc_13_00_1e_12_fc_11_15_11_00_f7_dd_f6_05_0d_f3_1a_13_fd_18_0e_f1_14_09_dd_0a_00_00_00_00_00_00_00_00_ed_e6_f1_06_ed_fc_fb_fe_10_07_f0_17_15_03_07_f5_0a_13_06_13_fa_1c_07_05_03_ee_eb_f1_00_00_00_00_00_00_00_00_dc_09_f6_fc_fb_04_d9_f9_08_01_08_18_15_25_e6_fe_f9_03_f1_fc_f3_fb_0e_00_f2_f0_0a_f7_00_00_00_00_00_00_00_00_06_0b_f8_26_f5_0c_e6_09_f7_fe_fa_04_fa_0b_dc_f8_12_e4_f3_f5_02_0a_f9_20_fd_04_12_fa_00_00_00_00_00_00_00_00_fb_03_15_e2_ef_f4_01_19_0c_fd_fc_fc_03_0f_18_f2_05_e9_f2_22_04_ef_f5_03_fd_10_f4_e2_00_00_00_00_00_00_00_00_0b_07_02_ec_f8_01_0e_fe_fc_03_ef_eb_f1_f9_04_06_09_15_fc_01_03_f9_0d_ec_f2_2a_e9_01_00_00_00_00_00_00_00_00_0b_12_e9_ff_e9_0d_f3_0f_e4_02_08_0d_e9_e3_fc_05_f3_f6_fd_ee_fc_e4_f5_f3_ef_e1_06_f5_00_00_00_00_00_00_00_00_0b_00_16_e1_f2_f1_06_03_ff_fa_07_f3_09_f7_0a_0a_0c_ff_1f_f4_0f_ef_fb_15_02_e6_fd_f9_00_00_00_00_00_00_00_00_08_f1_ff_f1_eb_11_f4_ea_fd_f3_f0_05_0a_e9_05_0a_f7_e8_f7_f2_11_f4_03_f5_13_e9_fb_fc_00_00_00_00_00_00_00_00_04_fb_0a_01_f9_04_00_03_f7_fb_0b_2c_13_0a_10_ec_08_eb_17_fa_1e_05_18_f4_02_01_0a_03_00_00_00_00_00_00_00_00_ff_02_f6_f9_f6_00_07_01_01_f2_0d_19_fc_05_ef_f3_0c_e7_0d_e1_07_09_26_ff_f8_0a_cf_f1_00_00_00_00_00_00_00_00_e9_08_04_ff_fe_e4_dc_fa_05_fc_23_09_ff_03_09_04_18_1a_f4_02_d7_2a_ed_09_07_14_f0_ff_00_00_00_00_00_00_00_00_0f_09_0f_f8_08_f1_21_02_27_fc_f8_fb_ef_11_ee_f9_17_13_01_2c_04_f6_1c_e8_f7_f8_fa_08_00_00_00_00_00_00_00_00_13_f6_11_24_fb_00_f4_09_0d_ff_ff_2c_f2_0f_2b_e0_fa_0c_04_25_fa_0a_0c_0c_15_f9_07_f6_00_00_00_00_00_00_00_00_fa_f7_07_20_f8_17_10_07_0a_07_1a_04_0b_f6_ff_1a_ef_e6_03_02_06_1f_fb_0c_06_f9_ff_04_00_00_00_00_00_00_00_00_1c_ec_f8_09_fc_20_e8_0e_f6_ed_f6_1c_00_e9_f6_07_15_f1_06_12_f9_e7_ef_08_ed_fb_16_fd_00_00_00_00_00_00_00_00_13_0d_fa_df_f0_09_e6_fd_f5_09_03_fa_17_fa_2f_16_ff_09_10_04_09_fe_fd_0d_f6_f2_e3_e2_00_00_00_00_00_00_00_00_f1_12_1b_ed_fb_18_fe_fd_01_1b_01_01_f3_1d_ff_07_0f_fe_05_ef_ef_38_fc_fb_ee_fc_f0_0e_00_00_00_00_00_00_00_00_02_37_0c_f4_1e_e1_04_f4_f4_0a_22_06_01_f0_00_00_1d_0d_fd_1f_f4_06_02_fe_07_ec_12_f7_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;

wire out_valid;
wire [image_size*image_size*word_length-1 :0] data_out;
wire [image_size*image_size*col_length-1:0] data_out_cols;
wire [image_size*image_size*col_length-1:0] data_out_rows;

wire [word_length-1:0] pixels_0_0, pixels_0_1, pixels_0_2, pixels_0_3, pixels_0_4, pixels_0_5, pixels_0_6, pixels_0_7, pixels_0_8, pixels_0_9, pixels_0_10, pixels_0_11, pixels_0_12, pixels_0_13, pixels_0_14, pixels_0_15, pixels_0_16, pixels_0_17, pixels_0_18, pixels_0_19, pixels_0_20, pixels_0_21, pixels_0_22, pixels_0_23, pixels_0_24, pixels_0_25, pixels_0_26, pixels_0_27, pixels_0_28, pixels_0_29, pixels_0_30, pixels_0_31, pixels_0_32, pixels_0_33, pixels_0_34, pixels_0_35, pixels_1_0, pixels_1_1, pixels_1_2, pixels_1_3, pixels_1_4, pixels_1_5, pixels_1_6, pixels_1_7, pixels_1_8, pixels_1_9, pixels_1_10, pixels_1_11, pixels_1_12, pixels_1_13, pixels_1_14, pixels_1_15, pixels_1_16, pixels_1_17, pixels_1_18, pixels_1_19, pixels_1_20, pixels_1_21, pixels_1_22, pixels_1_23, pixels_1_24, pixels_1_25, pixels_1_26, pixels_1_27, pixels_1_28, pixels_1_29, pixels_1_30, pixels_1_31, pixels_1_32, pixels_1_33, pixels_1_34, pixels_1_35, pixels_2_0, pixels_2_1, pixels_2_2, pixels_2_3, pixels_2_4, pixels_2_5, pixels_2_6, pixels_2_7, pixels_2_8, pixels_2_9, pixels_2_10, pixels_2_11, pixels_2_12, pixels_2_13, pixels_2_14, pixels_2_15, pixels_2_16, pixels_2_17, pixels_2_18, pixels_2_19, pixels_2_20, pixels_2_21, pixels_2_22, pixels_2_23, pixels_2_24, pixels_2_25, pixels_2_26, pixels_2_27, pixels_2_28, pixels_2_29, pixels_2_30, pixels_2_31, pixels_2_32, pixels_2_33, pixels_2_34, pixels_2_35, pixels_3_0, pixels_3_1, pixels_3_2, pixels_3_3, pixels_3_4, pixels_3_5, pixels_3_6, pixels_3_7, pixels_3_8, pixels_3_9, pixels_3_10, pixels_3_11, pixels_3_12, pixels_3_13, pixels_3_14, pixels_3_15, pixels_3_16, pixels_3_17, pixels_3_18, pixels_3_19, pixels_3_20, pixels_3_21, pixels_3_22, pixels_3_23, pixels_3_24, pixels_3_25, pixels_3_26, pixels_3_27, pixels_3_28, pixels_3_29, pixels_3_30, pixels_3_31, pixels_3_32, pixels_3_33, pixels_3_34, pixels_3_35, pixels_4_0, pixels_4_1, pixels_4_2, pixels_4_3, pixels_4_4, pixels_4_5, pixels_4_6, pixels_4_7, pixels_4_8, pixels_4_9, pixels_4_10, pixels_4_11, pixels_4_12, pixels_4_13, pixels_4_14, pixels_4_15, pixels_4_16, pixels_4_17, pixels_4_18, pixels_4_19, pixels_4_20, pixels_4_21, pixels_4_22, pixels_4_23, pixels_4_24, pixels_4_25, pixels_4_26, pixels_4_27, pixels_4_28, pixels_4_29, pixels_4_30, pixels_4_31, pixels_4_32, pixels_4_33, pixels_4_34, pixels_4_35, pixels_5_0, pixels_5_1, pixels_5_2, pixels_5_3, pixels_5_4, pixels_5_5, pixels_5_6, pixels_5_7, pixels_5_8, pixels_5_9, pixels_5_10, pixels_5_11, pixels_5_12, pixels_5_13, pixels_5_14, pixels_5_15, pixels_5_16, pixels_5_17, pixels_5_18, pixels_5_19, pixels_5_20, pixels_5_21, pixels_5_22, pixels_5_23, pixels_5_24, pixels_5_25, pixels_5_26, pixels_5_27, pixels_5_28, pixels_5_29, pixels_5_30, pixels_5_31, pixels_5_32, pixels_5_33, pixels_5_34, pixels_5_35, pixels_6_0, pixels_6_1, pixels_6_2, pixels_6_3, pixels_6_4, pixels_6_5, pixels_6_6, pixels_6_7, pixels_6_8, pixels_6_9, pixels_6_10, pixels_6_11, pixels_6_12, pixels_6_13, pixels_6_14, pixels_6_15, pixels_6_16, pixels_6_17, pixels_6_18, pixels_6_19, pixels_6_20, pixels_6_21, pixels_6_22, pixels_6_23, pixels_6_24, pixels_6_25, pixels_6_26, pixels_6_27, pixels_6_28, pixels_6_29, pixels_6_30, pixels_6_31, pixels_6_32, pixels_6_33, pixels_6_34, pixels_6_35, pixels_7_0, pixels_7_1, pixels_7_2, pixels_7_3, pixels_7_4, pixels_7_5, pixels_7_6, pixels_7_7, pixels_7_8, pixels_7_9, pixels_7_10, pixels_7_11, pixels_7_12, pixels_7_13, pixels_7_14, pixels_7_15, pixels_7_16, pixels_7_17, pixels_7_18, pixels_7_19, pixels_7_20, pixels_7_21, pixels_7_22, pixels_7_23, pixels_7_24, pixels_7_25, pixels_7_26, pixels_7_27, pixels_7_28, pixels_7_29, pixels_7_30, pixels_7_31, pixels_7_32, pixels_7_33, pixels_7_34, pixels_7_35, pixels_8_0, pixels_8_1, pixels_8_2, pixels_8_3, pixels_8_4, pixels_8_5, pixels_8_6, pixels_8_7, pixels_8_8, pixels_8_9, pixels_8_10, pixels_8_11, pixels_8_12, pixels_8_13, pixels_8_14, pixels_8_15, pixels_8_16, pixels_8_17, pixels_8_18, pixels_8_19, pixels_8_20, pixels_8_21, pixels_8_22, pixels_8_23, pixels_8_24, pixels_8_25, pixels_8_26, pixels_8_27, pixels_8_28, pixels_8_29, pixels_8_30, pixels_8_31, pixels_8_32, pixels_8_33, pixels_8_34, pixels_8_35, pixels_9_0, pixels_9_1, pixels_9_2, pixels_9_3, pixels_9_4, pixels_9_5, pixels_9_6, pixels_9_7, pixels_9_8, pixels_9_9, pixels_9_10, pixels_9_11, pixels_9_12, pixels_9_13, pixels_9_14, pixels_9_15, pixels_9_16, pixels_9_17, pixels_9_18, pixels_9_19, pixels_9_20, pixels_9_21, pixels_9_22, pixels_9_23, pixels_9_24, pixels_9_25, pixels_9_26, pixels_9_27, pixels_9_28, pixels_9_29, pixels_9_30, pixels_9_31, pixels_9_32, pixels_9_33, pixels_9_34, pixels_9_35, pixels_10_0, pixels_10_1, pixels_10_2, pixels_10_3, pixels_10_4, pixels_10_5, pixels_10_6, pixels_10_7, pixels_10_8, pixels_10_9, pixels_10_10, pixels_10_11, pixels_10_12, pixels_10_13, pixels_10_14, pixels_10_15, pixels_10_16, pixels_10_17, pixels_10_18, pixels_10_19, pixels_10_20, pixels_10_21, pixels_10_22, pixels_10_23, pixels_10_24, pixels_10_25, pixels_10_26, pixels_10_27, pixels_10_28, pixels_10_29, pixels_10_30, pixels_10_31, pixels_10_32, pixels_10_33, pixels_10_34, pixels_10_35, pixels_11_0, pixels_11_1, pixels_11_2, pixels_11_3, pixels_11_4, pixels_11_5, pixels_11_6, pixels_11_7, pixels_11_8, pixels_11_9, pixels_11_10, pixels_11_11, pixels_11_12, pixels_11_13, pixels_11_14, pixels_11_15, pixels_11_16, pixels_11_17, pixels_11_18, pixels_11_19, pixels_11_20, pixels_11_21, pixels_11_22, pixels_11_23, pixels_11_24, pixels_11_25, pixels_11_26, pixels_11_27, pixels_11_28, pixels_11_29, pixels_11_30, pixels_11_31, pixels_11_32, pixels_11_33, pixels_11_34, pixels_11_35, pixels_12_0, pixels_12_1, pixels_12_2, pixels_12_3, pixels_12_4, pixels_12_5, pixels_12_6, pixels_12_7, pixels_12_8, pixels_12_9, pixels_12_10, pixels_12_11, pixels_12_12, pixels_12_13, pixels_12_14, pixels_12_15, pixels_12_16, pixels_12_17, pixels_12_18, pixels_12_19, pixels_12_20, pixels_12_21, pixels_12_22, pixels_12_23, pixels_12_24, pixels_12_25, pixels_12_26, pixels_12_27, pixels_12_28, pixels_12_29, pixels_12_30, pixels_12_31, pixels_12_32, pixels_12_33, pixels_12_34, pixels_12_35, pixels_13_0, pixels_13_1, pixels_13_2, pixels_13_3, pixels_13_4, pixels_13_5, pixels_13_6, pixels_13_7, pixels_13_8, pixels_13_9, pixels_13_10, pixels_13_11, pixels_13_12, pixels_13_13, pixels_13_14, pixels_13_15, pixels_13_16, pixels_13_17, pixels_13_18, pixels_13_19, pixels_13_20, pixels_13_21, pixels_13_22, pixels_13_23, pixels_13_24, pixels_13_25, pixels_13_26, pixels_13_27, pixels_13_28, pixels_13_29, pixels_13_30, pixels_13_31, pixels_13_32, pixels_13_33, pixels_13_34, pixels_13_35, pixels_14_0, pixels_14_1, pixels_14_2, pixels_14_3, pixels_14_4, pixels_14_5, pixels_14_6, pixels_14_7, pixels_14_8, pixels_14_9, pixels_14_10, pixels_14_11, pixels_14_12, pixels_14_13, pixels_14_14, pixels_14_15, pixels_14_16, pixels_14_17, pixels_14_18, pixels_14_19, pixels_14_20, pixels_14_21, pixels_14_22, pixels_14_23, pixels_14_24, pixels_14_25, pixels_14_26, pixels_14_27, pixels_14_28, pixels_14_29, pixels_14_30, pixels_14_31, pixels_14_32, pixels_14_33, pixels_14_34, pixels_14_35, pixels_15_0, pixels_15_1, pixels_15_2, pixels_15_3, pixels_15_4, pixels_15_5, pixels_15_6, pixels_15_7, pixels_15_8, pixels_15_9, pixels_15_10, pixels_15_11, pixels_15_12, pixels_15_13, pixels_15_14, pixels_15_15, pixels_15_16, pixels_15_17, pixels_15_18, pixels_15_19, pixels_15_20, pixels_15_21, pixels_15_22, pixels_15_23, pixels_15_24, pixels_15_25, pixels_15_26, pixels_15_27, pixels_15_28, pixels_15_29, pixels_15_30, pixels_15_31, pixels_15_32, pixels_15_33, pixels_15_34, pixels_15_35, pixels_16_0, pixels_16_1, pixels_16_2, pixels_16_3, pixels_16_4, pixels_16_5, pixels_16_6, pixels_16_7, pixels_16_8, pixels_16_9, pixels_16_10, pixels_16_11, pixels_16_12, pixels_16_13, pixels_16_14, pixels_16_15, pixels_16_16, pixels_16_17, pixels_16_18, pixels_16_19, pixels_16_20, pixels_16_21, pixels_16_22, pixels_16_23, pixels_16_24, pixels_16_25, pixels_16_26, pixels_16_27, pixels_16_28, pixels_16_29, pixels_16_30, pixels_16_31, pixels_16_32, pixels_16_33, pixels_16_34, pixels_16_35, pixels_17_0, pixels_17_1, pixels_17_2, pixels_17_3, pixels_17_4, pixels_17_5, pixels_17_6, pixels_17_7, pixels_17_8, pixels_17_9, pixels_17_10, pixels_17_11, pixels_17_12, pixels_17_13, pixels_17_14, pixels_17_15, pixels_17_16, pixels_17_17, pixels_17_18, pixels_17_19, pixels_17_20, pixels_17_21, pixels_17_22, pixels_17_23, pixels_17_24, pixels_17_25, pixels_17_26, pixels_17_27, pixels_17_28, pixels_17_29, pixels_17_30, pixels_17_31, pixels_17_32, pixels_17_33, pixels_17_34, pixels_17_35, pixels_18_0, pixels_18_1, pixels_18_2, pixels_18_3, pixels_18_4, pixels_18_5, pixels_18_6, pixels_18_7, pixels_18_8, pixels_18_9, pixels_18_10, pixels_18_11, pixels_18_12, pixels_18_13, pixels_18_14, pixels_18_15, pixels_18_16, pixels_18_17, pixels_18_18, pixels_18_19, pixels_18_20, pixels_18_21, pixels_18_22, pixels_18_23, pixels_18_24, pixels_18_25, pixels_18_26, pixels_18_27, pixels_18_28, pixels_18_29, pixels_18_30, pixels_18_31, pixels_18_32, pixels_18_33, pixels_18_34, pixels_18_35, pixels_19_0, pixels_19_1, pixels_19_2, pixels_19_3, pixels_19_4, pixels_19_5, pixels_19_6, pixels_19_7, pixels_19_8, pixels_19_9, pixels_19_10, pixels_19_11, pixels_19_12, pixels_19_13, pixels_19_14, pixels_19_15, pixels_19_16, pixels_19_17, pixels_19_18, pixels_19_19, pixels_19_20, pixels_19_21, pixels_19_22, pixels_19_23, pixels_19_24, pixels_19_25, pixels_19_26, pixels_19_27, pixels_19_28, pixels_19_29, pixels_19_30, pixels_19_31, pixels_19_32, pixels_19_33, pixels_19_34, pixels_19_35, pixels_20_0, pixels_20_1, pixels_20_2, pixels_20_3, pixels_20_4, pixels_20_5, pixels_20_6, pixels_20_7, pixels_20_8, pixels_20_9, pixels_20_10, pixels_20_11, pixels_20_12, pixels_20_13, pixels_20_14, pixels_20_15, pixels_20_16, pixels_20_17, pixels_20_18, pixels_20_19, pixels_20_20, pixels_20_21, pixels_20_22, pixels_20_23, pixels_20_24, pixels_20_25, pixels_20_26, pixels_20_27, pixels_20_28, pixels_20_29, pixels_20_30, pixels_20_31, 
pixels_20_32, pixels_20_33, pixels_20_34, pixels_20_35, pixels_21_0, pixels_21_1, pixels_21_2, pixels_21_3, pixels_21_4, pixels_21_5, pixels_21_6, pixels_21_7, pixels_21_8, pixels_21_9, pixels_21_10, pixels_21_11, pixels_21_12, pixels_21_13, pixels_21_14, pixels_21_15, pixels_21_16, pixels_21_17, pixels_21_18, pixels_21_19, pixels_21_20, pixels_21_21, pixels_21_22, pixels_21_23, pixels_21_24, pixels_21_25, pixels_21_26, pixels_21_27, pixels_21_28, pixels_21_29, pixels_21_30, pixels_21_31, pixels_21_32, pixels_21_33, pixels_21_34, pixels_21_35, pixels_22_0, pixels_22_1, pixels_22_2, pixels_22_3, pixels_22_4, pixels_22_5, pixels_22_6, pixels_22_7, pixels_22_8, pixels_22_9, pixels_22_10, pixels_22_11, pixels_22_12, pixels_22_13, pixels_22_14, pixels_22_15, pixels_22_16, pixels_22_17, pixels_22_18, pixels_22_19, pixels_22_20, pixels_22_21, pixels_22_22, pixels_22_23, pixels_22_24, pixels_22_25, pixels_22_26, pixels_22_27, pixels_22_28, pixels_22_29, pixels_22_30, pixels_22_31, pixels_22_32, pixels_22_33, pixels_22_34, pixels_22_35, pixels_23_0, pixels_23_1, pixels_23_2, pixels_23_3, pixels_23_4, pixels_23_5, pixels_23_6, pixels_23_7, pixels_23_8, pixels_23_9, pixels_23_10, pixels_23_11, pixels_23_12, pixels_23_13, pixels_23_14, pixels_23_15, pixels_23_16, pixels_23_17, pixels_23_18, pixels_23_19, pixels_23_20, pixels_23_21, pixels_23_22, pixels_23_23, pixels_23_24, pixels_23_25, pixels_23_26, pixels_23_27, pixels_23_28, pixels_23_29, pixels_23_30, pixels_23_31, pixels_23_32, pixels_23_33, pixels_23_34, pixels_23_35, pixels_24_0, pixels_24_1, pixels_24_2, pixels_24_3, pixels_24_4, pixels_24_5, pixels_24_6, pixels_24_7, pixels_24_8, pixels_24_9, pixels_24_10, pixels_24_11, pixels_24_12, pixels_24_13, pixels_24_14, pixels_24_15, pixels_24_16, pixels_24_17, pixels_24_18, pixels_24_19, pixels_24_20, pixels_24_21, pixels_24_22, pixels_24_23, pixels_24_24, pixels_24_25, pixels_24_26, pixels_24_27, pixels_24_28, pixels_24_29, pixels_24_30, pixels_24_31, pixels_24_32, pixels_24_33, pixels_24_34, pixels_24_35, pixels_25_0, pixels_25_1, pixels_25_2, pixels_25_3, pixels_25_4, pixels_25_5, pixels_25_6, pixels_25_7, pixels_25_8, pixels_25_9, pixels_25_10, pixels_25_11, pixels_25_12, pixels_25_13, pixels_25_14, pixels_25_15, pixels_25_16, pixels_25_17, pixels_25_18, pixels_25_19, pixels_25_20, pixels_25_21, pixels_25_22, pixels_25_23, pixels_25_24, pixels_25_25, pixels_25_26, pixels_25_27, pixels_25_28, pixels_25_29, pixels_25_30, pixels_25_31, pixels_25_32, pixels_25_33, pixels_25_34, pixels_25_35, pixels_26_0, pixels_26_1, pixels_26_2, pixels_26_3, pixels_26_4, pixels_26_5, pixels_26_6, pixels_26_7, pixels_26_8, pixels_26_9, pixels_26_10, pixels_26_11, pixels_26_12, pixels_26_13, pixels_26_14, pixels_26_15, pixels_26_16, pixels_26_17, pixels_26_18, pixels_26_19, pixels_26_20, pixels_26_21, pixels_26_22, pixels_26_23, pixels_26_24, pixels_26_25, pixels_26_26, pixels_26_27, pixels_26_28, pixels_26_29, pixels_26_30, pixels_26_31, pixels_26_32, pixels_26_33, pixels_26_34, pixels_26_35, pixels_27_0, pixels_27_1, pixels_27_2, pixels_27_3, pixels_27_4, pixels_27_5, pixels_27_6, pixels_27_7, pixels_27_8, pixels_27_9, pixels_27_10, pixels_27_11, pixels_27_12, pixels_27_13, pixels_27_14, pixels_27_15, pixels_27_16, pixels_27_17, pixels_27_18, pixels_27_19, pixels_27_20, pixels_27_21, pixels_27_22, pixels_27_23, pixels_27_24, pixels_27_25, pixels_27_26, pixels_27_27, pixels_27_28, pixels_27_29, pixels_27_30, pixels_27_31, pixels_27_32, pixels_27_33, pixels_27_34, pixels_27_35, pixels_28_0, pixels_28_1, pixels_28_2, pixels_28_3, pixels_28_4, pixels_28_5, pixels_28_6, pixels_28_7, pixels_28_8, pixels_28_9, pixels_28_10, pixels_28_11, pixels_28_12, pixels_28_13, pixels_28_14, pixels_28_15, pixels_28_16, pixels_28_17, pixels_28_18, pixels_28_19, pixels_28_20, pixels_28_21, pixels_28_22, pixels_28_23, pixels_28_24, pixels_28_25, pixels_28_26, pixels_28_27, pixels_28_28, pixels_28_29, pixels_28_30, pixels_28_31, pixels_28_32, pixels_28_33, pixels_28_34, pixels_28_35, pixels_29_0, pixels_29_1, pixels_29_2, pixels_29_3, pixels_29_4, pixels_29_5, pixels_29_6, pixels_29_7, pixels_29_8, pixels_29_9, pixels_29_10, pixels_29_11, pixels_29_12, pixels_29_13, pixels_29_14, pixels_29_15, pixels_29_16, pixels_29_17, pixels_29_18, pixels_29_19, pixels_29_20, pixels_29_21, pixels_29_22, pixels_29_23, pixels_29_24, pixels_29_25, pixels_29_26, pixels_29_27, pixels_29_28, pixels_29_29, pixels_29_30, pixels_29_31, pixels_29_32, pixels_29_33, pixels_29_34, pixels_29_35, pixels_30_0, pixels_30_1, pixels_30_2, pixels_30_3, pixels_30_4, pixels_30_5, pixels_30_6, pixels_30_7, pixels_30_8, pixels_30_9, pixels_30_10, pixels_30_11, pixels_30_12, pixels_30_13, pixels_30_14, pixels_30_15, pixels_30_16, pixels_30_17, pixels_30_18, pixels_30_19, pixels_30_20, pixels_30_21, pixels_30_22, pixels_30_23, pixels_30_24, pixels_30_25, pixels_30_26, pixels_30_27, pixels_30_28, pixels_30_29, pixels_30_30, pixels_30_31, pixels_30_32, pixels_30_33, pixels_30_34, pixels_30_35, pixels_31_0, pixels_31_1, pixels_31_2, pixels_31_3, pixels_31_4, pixels_31_5, pixels_31_6, pixels_31_7, pixels_31_8, pixels_31_9, pixels_31_10, pixels_31_11, pixels_31_12, pixels_31_13, pixels_31_14, pixels_31_15, pixels_31_16, pixels_31_17, pixels_31_18, pixels_31_19, pixels_31_20, pixels_31_21, pixels_31_22, pixels_31_23, pixels_31_24, pixels_31_25, pixels_31_26, pixels_31_27, pixels_31_28, pixels_31_29, pixels_31_30, pixels_31_31, pixels_31_32, pixels_31_33, pixels_31_34, pixels_31_35, pixels_32_0, pixels_32_1, pixels_32_2, pixels_32_3, pixels_32_4, pixels_32_5, pixels_32_6, pixels_32_7, pixels_32_8, pixels_32_9, pixels_32_10, pixels_32_11, pixels_32_12, pixels_32_13, pixels_32_14, pixels_32_15, pixels_32_16, pixels_32_17, pixels_32_18, pixels_32_19, pixels_32_20, pixels_32_21, pixels_32_22, pixels_32_23, pixels_32_24, pixels_32_25, pixels_32_26, pixels_32_27, pixels_32_28, pixels_32_29, pixels_32_30, pixels_32_31, pixels_32_32, pixels_32_33, pixels_32_34, pixels_32_35, pixels_33_0, pixels_33_1, pixels_33_2, pixels_33_3, pixels_33_4, pixels_33_5, pixels_33_6, pixels_33_7, pixels_33_8, pixels_33_9, pixels_33_10, pixels_33_11, pixels_33_12, pixels_33_13, pixels_33_14, pixels_33_15, pixels_33_16, pixels_33_17, pixels_33_18, pixels_33_19, pixels_33_20, pixels_33_21, pixels_33_22, pixels_33_23, pixels_33_24, pixels_33_25, pixels_33_26, pixels_33_27, pixels_33_28, pixels_33_29, pixels_33_30, pixels_33_31, pixels_33_32, pixels_33_33, pixels_33_34, pixels_33_35, pixels_34_0, pixels_34_1, pixels_34_2, pixels_34_3, pixels_34_4, pixels_34_5, pixels_34_6, pixels_34_7, pixels_34_8, pixels_34_9, pixels_34_10, pixels_34_11, pixels_34_12, pixels_34_13, pixels_34_14, pixels_34_15, pixels_34_16, pixels_34_17, pixels_34_18, pixels_34_19, pixels_34_20, pixels_34_21, pixels_34_22, pixels_34_23, pixels_34_24, pixels_34_25, pixels_34_26, pixels_34_27, pixels_34_28, pixels_34_29, pixels_34_30, pixels_34_31, pixels_34_32, pixels_34_33, pixels_34_34, pixels_34_35, pixels_35_0, pixels_35_1, pixels_35_2, pixels_35_3, pixels_35_4, pixels_35_5, pixels_35_6, pixels_35_7, pixels_35_8, pixels_35_9, pixels_35_10, pixels_35_11, pixels_35_12, pixels_35_13, pixels_35_14, pixels_35_15, pixels_35_16, pixels_35_17, pixels_35_18, pixels_35_19, pixels_35_20, pixels_35_21, pixels_35_22, pixels_35_23, pixels_35_24, pixels_35_25, pixels_35_26, pixels_35_27, pixels_35_28, pixels_35_29, pixels_35_30, pixels_35_31, pixels_35_32, pixels_35_33, pixels_35_34, pixels_35_35;
assign pixels_0_0 = {data_out[1*word_length-1 -: word_length]};
assign pixels_0_1 = {data_out[2*word_length-1 -: word_length]};
assign pixels_0_2 = {data_out[3*word_length-1 -: word_length]};
assign pixels_0_3 = {data_out[4*word_length-1 -: word_length]};
assign pixels_0_4 = {data_out[5*word_length-1 -: word_length]};
assign pixels_0_5 = {data_out[6*word_length-1 -: word_length]};
assign pixels_0_6 = {data_out[7*word_length-1 -: word_length]};
assign pixels_0_7 = {data_out[8*word_length-1 -: word_length]};
assign pixels_0_8 = {data_out[9*word_length-1 -: word_length]};
assign pixels_0_9 = {data_out[10*word_length-1 -: word_length]};
assign pixels_0_10 = {data_out[11*word_length-1 -: word_length]};
assign pixels_0_11 = {data_out[12*word_length-1 -: word_length]};
assign pixels_0_12 = {data_out[13*word_length-1 -: word_length]};
assign pixels_0_13 = {data_out[14*word_length-1 -: word_length]};
assign pixels_0_14 = {data_out[15*word_length-1 -: word_length]};
assign pixels_0_15 = {data_out[16*word_length-1 -: word_length]};
assign pixels_0_16 = {data_out[17*word_length-1 -: word_length]};
assign pixels_0_17 = {data_out[18*word_length-1 -: word_length]};
assign pixels_0_18 = {data_out[19*word_length-1 -: word_length]};
assign pixels_0_19 = {data_out[20*word_length-1 -: word_length]};
assign pixels_0_20 = {data_out[21*word_length-1 -: word_length]};
assign pixels_0_21 = {data_out[22*word_length-1 -: word_length]};
assign pixels_0_22 = {data_out[23*word_length-1 -: word_length]};
assign pixels_0_23 = {data_out[24*word_length-1 -: word_length]};
assign pixels_0_24 = {data_out[25*word_length-1 -: word_length]};
assign pixels_0_25 = {data_out[26*word_length-1 -: word_length]};
assign pixels_0_26 = {data_out[27*word_length-1 -: word_length]};
assign pixels_0_27 = {data_out[28*word_length-1 -: word_length]};
assign pixels_0_28 = {data_out[29*word_length-1 -: word_length]};
assign pixels_0_29 = {data_out[30*word_length-1 -: word_length]};
assign pixels_0_30 = {data_out[31*word_length-1 -: word_length]};
assign pixels_0_31 = {data_out[32*word_length-1 -: word_length]};
assign pixels_0_32 = {data_out[33*word_length-1 -: word_length]};
assign pixels_0_33 = {data_out[34*word_length-1 -: word_length]};
assign pixels_0_34 = {data_out[35*word_length-1 -: word_length]};
assign pixels_0_35 = {data_out[36*word_length-1 -: word_length]};
assign pixels_1_0 = {data_out[37*word_length-1 -: word_length]};
assign pixels_1_1 = {data_out[38*word_length-1 -: word_length]};
assign pixels_1_2 = {data_out[39*word_length-1 -: word_length]};
assign pixels_1_3 = {data_out[40*word_length-1 -: word_length]};
assign pixels_1_4 = {data_out[41*word_length-1 -: word_length]};
assign pixels_1_5 = {data_out[42*word_length-1 -: word_length]};
assign pixels_1_6 = {data_out[43*word_length-1 -: word_length]};
assign pixels_1_7 = {data_out[44*word_length-1 -: word_length]};
assign pixels_1_8 = {data_out[45*word_length-1 -: word_length]};
assign pixels_1_9 = {data_out[46*word_length-1 -: word_length]};
assign pixels_1_10 = {data_out[47*word_length-1 -: word_length]};
assign pixels_1_11 = {data_out[48*word_length-1 -: word_length]};
assign pixels_1_12 = {data_out[49*word_length-1 -: word_length]};
assign pixels_1_13 = {data_out[50*word_length-1 -: word_length]};
assign pixels_1_14 = {data_out[51*word_length-1 -: word_length]};
assign pixels_1_15 = {data_out[52*word_length-1 -: word_length]};
assign pixels_1_16 = {data_out[53*word_length-1 -: word_length]};
assign pixels_1_17 = {data_out[54*word_length-1 -: word_length]};
assign pixels_1_18 = {data_out[55*word_length-1 -: word_length]};
assign pixels_1_19 = {data_out[56*word_length-1 -: word_length]};
assign pixels_1_20 = {data_out[57*word_length-1 -: word_length]};
assign pixels_1_21 = {data_out[58*word_length-1 -: word_length]};
assign pixels_1_22 = {data_out[59*word_length-1 -: word_length]};
assign pixels_1_23 = {data_out[60*word_length-1 -: word_length]};
assign pixels_1_24 = {data_out[61*word_length-1 -: word_length]};
assign pixels_1_25 = {data_out[62*word_length-1 -: word_length]};
assign pixels_1_26 = {data_out[63*word_length-1 -: word_length]};
assign pixels_1_27 = {data_out[64*word_length-1 -: word_length]};
assign pixels_1_28 = {data_out[65*word_length-1 -: word_length]};
assign pixels_1_29 = {data_out[66*word_length-1 -: word_length]};
assign pixels_1_30 = {data_out[67*word_length-1 -: word_length]};
assign pixels_1_31 = {data_out[68*word_length-1 -: word_length]};
assign pixels_1_32 = {data_out[69*word_length-1 -: word_length]};
assign pixels_1_33 = {data_out[70*word_length-1 -: word_length]};
assign pixels_1_34 = {data_out[71*word_length-1 -: word_length]};
assign pixels_1_35 = {data_out[72*word_length-1 -: word_length]};
assign pixels_2_0 = {data_out[73*word_length-1 -: word_length]};
assign pixels_2_1 = {data_out[74*word_length-1 -: word_length]};
assign pixels_2_2 = {data_out[75*word_length-1 -: word_length]};
assign pixels_2_3 = {data_out[76*word_length-1 -: word_length]};
assign pixels_2_4 = {data_out[77*word_length-1 -: word_length]};
assign pixels_2_5 = {data_out[78*word_length-1 -: word_length]};
assign pixels_2_6 = {data_out[79*word_length-1 -: word_length]};
assign pixels_2_7 = {data_out[80*word_length-1 -: word_length]};
assign pixels_2_8 = {data_out[81*word_length-1 -: word_length]};
assign pixels_2_9 = {data_out[82*word_length-1 -: word_length]};
assign pixels_2_10 = {data_out[83*word_length-1 -: word_length]};
assign pixels_2_11 = {data_out[84*word_length-1 -: word_length]};
assign pixels_2_12 = {data_out[85*word_length-1 -: word_length]};
assign pixels_2_13 = {data_out[86*word_length-1 -: word_length]};
assign pixels_2_14 = {data_out[87*word_length-1 -: word_length]};
assign pixels_2_15 = {data_out[88*word_length-1 -: word_length]};
assign pixels_2_16 = {data_out[89*word_length-1 -: word_length]};
assign pixels_2_17 = {data_out[90*word_length-1 -: word_length]};
assign pixels_2_18 = {data_out[91*word_length-1 -: word_length]};
assign pixels_2_19 = {data_out[92*word_length-1 -: word_length]};
assign pixels_2_20 = {data_out[93*word_length-1 -: word_length]};
assign pixels_2_21 = {data_out[94*word_length-1 -: word_length]};
assign pixels_2_22 = {data_out[95*word_length-1 -: word_length]};
assign pixels_2_23 = {data_out[96*word_length-1 -: word_length]};
assign pixels_2_24 = {data_out[97*word_length-1 -: word_length]};
assign pixels_2_25 = {data_out[98*word_length-1 -: word_length]};
assign pixels_2_26 = {data_out[99*word_length-1 -: word_length]};
assign pixels_2_27 = {data_out[100*word_length-1 -: word_length]};
assign pixels_2_28 = {data_out[101*word_length-1 -: word_length]};
assign pixels_2_29 = {data_out[102*word_length-1 -: word_length]};
assign pixels_2_30 = {data_out[103*word_length-1 -: word_length]};
assign pixels_2_31 = {data_out[104*word_length-1 -: word_length]};
assign pixels_2_32 = {data_out[105*word_length-1 -: word_length]};
assign pixels_2_33 = {data_out[106*word_length-1 -: word_length]};
assign pixels_2_34 = {data_out[107*word_length-1 -: word_length]};
assign pixels_2_35 = {data_out[108*word_length-1 -: word_length]};
assign pixels_3_0 = {data_out[109*word_length-1 -: word_length]};
assign pixels_3_1 = {data_out[110*word_length-1 -: word_length]};
assign pixels_3_2 = {data_out[111*word_length-1 -: word_length]};
assign pixels_3_3 = {data_out[112*word_length-1 -: word_length]};
assign pixels_3_4 = {data_out[113*word_length-1 -: word_length]};
assign pixels_3_5 = {data_out[114*word_length-1 -: word_length]};
assign pixels_3_6 = {data_out[115*word_length-1 -: word_length]};
assign pixels_3_7 = {data_out[116*word_length-1 -: word_length]};
assign pixels_3_8 = {data_out[117*word_length-1 -: word_length]};
assign pixels_3_9 = {data_out[118*word_length-1 -: word_length]};
assign pixels_3_10 = {data_out[119*word_length-1 -: word_length]};
assign pixels_3_11 = {data_out[120*word_length-1 -: word_length]};
assign pixels_3_12 = {data_out[121*word_length-1 -: word_length]};
assign pixels_3_13 = {data_out[122*word_length-1 -: word_length]};
assign pixels_3_14 = {data_out[123*word_length-1 -: word_length]};
assign pixels_3_15 = {data_out[124*word_length-1 -: word_length]};
assign pixels_3_16 = {data_out[125*word_length-1 -: word_length]};
assign pixels_3_17 = {data_out[126*word_length-1 -: word_length]};
assign pixels_3_18 = {data_out[127*word_length-1 -: word_length]};
assign pixels_3_19 = {data_out[128*word_length-1 -: word_length]};
assign pixels_3_20 = {data_out[129*word_length-1 -: word_length]};
assign pixels_3_21 = {data_out[130*word_length-1 -: word_length]};
assign pixels_3_22 = {data_out[131*word_length-1 -: word_length]};
assign pixels_3_23 = {data_out[132*word_length-1 -: word_length]};
assign pixels_3_24 = {data_out[133*word_length-1 -: word_length]};
assign pixels_3_25 = {data_out[134*word_length-1 -: word_length]};
assign pixels_3_26 = {data_out[135*word_length-1 -: word_length]};
assign pixels_3_27 = {data_out[136*word_length-1 -: word_length]};
assign pixels_3_28 = {data_out[137*word_length-1 -: word_length]};
assign pixels_3_29 = {data_out[138*word_length-1 -: word_length]};
assign pixels_3_30 = {data_out[139*word_length-1 -: word_length]};
assign pixels_3_31 = {data_out[140*word_length-1 -: word_length]};
assign pixels_3_32 = {data_out[141*word_length-1 -: word_length]};
assign pixels_3_33 = {data_out[142*word_length-1 -: word_length]};
assign pixels_3_34 = {data_out[143*word_length-1 -: word_length]};
assign pixels_3_35 = {data_out[144*word_length-1 -: word_length]};
assign pixels_4_0 = {data_out[145*word_length-1 -: word_length]};
assign pixels_4_1 = {data_out[146*word_length-1 -: word_length]};
assign pixels_4_2 = {data_out[147*word_length-1 -: word_length]};
assign pixels_4_3 = {data_out[148*word_length-1 -: word_length]};
assign pixels_4_4 = {data_out[149*word_length-1 -: word_length]};
assign pixels_4_5 = {data_out[150*word_length-1 -: word_length]};
assign pixels_4_6 = {data_out[151*word_length-1 -: word_length]};
assign pixels_4_7 = {data_out[152*word_length-1 -: word_length]};
assign pixels_4_8 = {data_out[153*word_length-1 -: word_length]};
assign pixels_4_9 = {data_out[154*word_length-1 -: word_length]};
assign pixels_4_10 = {data_out[155*word_length-1 -: word_length]};
assign pixels_4_11 = {data_out[156*word_length-1 -: word_length]};
assign pixels_4_12 = {data_out[157*word_length-1 -: word_length]};
assign pixels_4_13 = {data_out[158*word_length-1 -: word_length]};
assign pixels_4_14 = {data_out[159*word_length-1 -: word_length]};
assign pixels_4_15 = {data_out[160*word_length-1 -: word_length]};
assign pixels_4_16 = {data_out[161*word_length-1 -: word_length]};
assign pixels_4_17 = {data_out[162*word_length-1 -: word_length]};
assign pixels_4_18 = {data_out[163*word_length-1 -: word_length]};
assign pixels_4_19 = {data_out[164*word_length-1 -: word_length]};
assign pixels_4_20 = {data_out[165*word_length-1 -: word_length]};
assign pixels_4_21 = {data_out[166*word_length-1 -: word_length]};
assign pixels_4_22 = {data_out[167*word_length-1 -: word_length]};
assign pixels_4_23 = {data_out[168*word_length-1 -: word_length]};
assign pixels_4_24 = {data_out[169*word_length-1 -: word_length]};
assign pixels_4_25 = {data_out[170*word_length-1 -: word_length]};
assign pixels_4_26 = {data_out[171*word_length-1 -: word_length]};
assign pixels_4_27 = {data_out[172*word_length-1 -: word_length]};
assign pixels_4_28 = {data_out[173*word_length-1 -: word_length]};
assign pixels_4_29 = {data_out[174*word_length-1 -: word_length]};
assign pixels_4_30 = {data_out[175*word_length-1 -: word_length]};
assign pixels_4_31 = {data_out[176*word_length-1 -: word_length]};
assign pixels_4_32 = {data_out[177*word_length-1 -: word_length]};
assign pixels_4_33 = {data_out[178*word_length-1 -: word_length]};
assign pixels_4_34 = {data_out[179*word_length-1 -: word_length]};
assign pixels_4_35 = {data_out[180*word_length-1 -: word_length]};
assign pixels_5_0 = {data_out[181*word_length-1 -: word_length]};
assign pixels_5_1 = {data_out[182*word_length-1 -: word_length]};
assign pixels_5_2 = {data_out[183*word_length-1 -: word_length]};
assign pixels_5_3 = {data_out[184*word_length-1 -: word_length]};
assign pixels_5_4 = {data_out[185*word_length-1 -: word_length]};
assign pixels_5_5 = {data_out[186*word_length-1 -: word_length]};
assign pixels_5_6 = {data_out[187*word_length-1 -: word_length]};
assign pixels_5_7 = {data_out[188*word_length-1 -: word_length]};
assign pixels_5_8 = {data_out[189*word_length-1 -: word_length]};
assign pixels_5_9 = {data_out[190*word_length-1 -: word_length]};
assign pixels_5_10 = {data_out[191*word_length-1 -: word_length]};
assign pixels_5_11 = {data_out[192*word_length-1 -: word_length]};
assign pixels_5_12 = {data_out[193*word_length-1 -: word_length]};
assign pixels_5_13 = {data_out[194*word_length-1 -: word_length]};
assign pixels_5_14 = {data_out[195*word_length-1 -: word_length]};
assign pixels_5_15 = {data_out[196*word_length-1 -: word_length]};
assign pixels_5_16 = {data_out[197*word_length-1 -: word_length]};
assign pixels_5_17 = {data_out[198*word_length-1 -: word_length]};
assign pixels_5_18 = {data_out[199*word_length-1 -: word_length]};
assign pixels_5_19 = {data_out[200*word_length-1 -: word_length]};
assign pixels_5_20 = {data_out[201*word_length-1 -: word_length]};
assign pixels_5_21 = {data_out[202*word_length-1 -: word_length]};
assign pixels_5_22 = {data_out[203*word_length-1 -: word_length]};
assign pixels_5_23 = {data_out[204*word_length-1 -: word_length]};
assign pixels_5_24 = {data_out[205*word_length-1 -: word_length]};
assign pixels_5_25 = {data_out[206*word_length-1 -: word_length]};
assign pixels_5_26 = {data_out[207*word_length-1 -: word_length]};
assign pixels_5_27 = {data_out[208*word_length-1 -: word_length]};
assign pixels_5_28 = {data_out[209*word_length-1 -: word_length]};
assign pixels_5_29 = {data_out[210*word_length-1 -: word_length]};
assign pixels_5_30 = {data_out[211*word_length-1 -: word_length]};
assign pixels_5_31 = {data_out[212*word_length-1 -: word_length]};
assign pixels_5_32 = {data_out[213*word_length-1 -: word_length]};
assign pixels_5_33 = {data_out[214*word_length-1 -: word_length]};
assign pixels_5_34 = {data_out[215*word_length-1 -: word_length]};
assign pixels_5_35 = {data_out[216*word_length-1 -: word_length]};
assign pixels_6_0 = {data_out[217*word_length-1 -: word_length]};
assign pixels_6_1 = {data_out[218*word_length-1 -: word_length]};
assign pixels_6_2 = {data_out[219*word_length-1 -: word_length]};
assign pixels_6_3 = {data_out[220*word_length-1 -: word_length]};
assign pixels_6_4 = {data_out[221*word_length-1 -: word_length]};
assign pixels_6_5 = {data_out[222*word_length-1 -: word_length]};
assign pixels_6_6 = {data_out[223*word_length-1 -: word_length]};
assign pixels_6_7 = {data_out[224*word_length-1 -: word_length]};
assign pixels_6_8 = {data_out[225*word_length-1 -: word_length]};
assign pixels_6_9 = {data_out[226*word_length-1 -: word_length]};
assign pixels_6_10 = {data_out[227*word_length-1 -: word_length]};
assign pixels_6_11 = {data_out[228*word_length-1 -: word_length]};
assign pixels_6_12 = {data_out[229*word_length-1 -: word_length]};
assign pixels_6_13 = {data_out[230*word_length-1 -: word_length]};
assign pixels_6_14 = {data_out[231*word_length-1 -: word_length]};
assign pixels_6_15 = {data_out[232*word_length-1 -: word_length]};
assign pixels_6_16 = {data_out[233*word_length-1 -: word_length]};
assign pixels_6_17 = {data_out[234*word_length-1 -: word_length]};
assign pixels_6_18 = {data_out[235*word_length-1 -: word_length]};
assign pixels_6_19 = {data_out[236*word_length-1 -: word_length]};
assign pixels_6_20 = {data_out[237*word_length-1 -: word_length]};
assign pixels_6_21 = {data_out[238*word_length-1 -: word_length]};
assign pixels_6_22 = {data_out[239*word_length-1 -: word_length]};
assign pixels_6_23 = {data_out[240*word_length-1 -: word_length]};
assign pixels_6_24 = {data_out[241*word_length-1 -: word_length]};
assign pixels_6_25 = {data_out[242*word_length-1 -: word_length]};
assign pixels_6_26 = {data_out[243*word_length-1 -: word_length]};
assign pixels_6_27 = {data_out[244*word_length-1 -: word_length]};
assign pixels_6_28 = {data_out[245*word_length-1 -: word_length]};
assign pixels_6_29 = {data_out[246*word_length-1 -: word_length]};
assign pixels_6_30 = {data_out[247*word_length-1 -: word_length]};
assign pixels_6_31 = {data_out[248*word_length-1 -: word_length]};
assign pixels_6_32 = {data_out[249*word_length-1 -: word_length]};
assign pixels_6_33 = {data_out[250*word_length-1 -: word_length]};
assign pixels_6_34 = {data_out[251*word_length-1 -: word_length]};
assign pixels_6_35 = {data_out[252*word_length-1 -: word_length]};
assign pixels_7_0 = {data_out[253*word_length-1 -: word_length]};
assign pixels_7_1 = {data_out[254*word_length-1 -: word_length]};
assign pixels_7_2 = {data_out[255*word_length-1 -: word_length]};
assign pixels_7_3 = {data_out[256*word_length-1 -: word_length]};
assign pixels_7_4 = {data_out[257*word_length-1 -: word_length]};
assign pixels_7_5 = {data_out[258*word_length-1 -: word_length]};
assign pixels_7_6 = {data_out[259*word_length-1 -: word_length]};
assign pixels_7_7 = {data_out[260*word_length-1 -: word_length]};
assign pixels_7_8 = {data_out[261*word_length-1 -: word_length]};
assign pixels_7_9 = {data_out[262*word_length-1 -: word_length]};
assign pixels_7_10 = {data_out[263*word_length-1 -: word_length]};
assign pixels_7_11 = {data_out[264*word_length-1 -: word_length]};
assign pixels_7_12 = {data_out[265*word_length-1 -: word_length]};
assign pixels_7_13 = {data_out[266*word_length-1 -: word_length]};
assign pixels_7_14 = {data_out[267*word_length-1 -: word_length]};
assign pixels_7_15 = {data_out[268*word_length-1 -: word_length]};
assign pixels_7_16 = {data_out[269*word_length-1 -: word_length]};
assign pixels_7_17 = {data_out[270*word_length-1 -: word_length]};
assign pixels_7_18 = {data_out[271*word_length-1 -: word_length]};
assign pixels_7_19 = {data_out[272*word_length-1 -: word_length]};
assign pixels_7_20 = {data_out[273*word_length-1 -: word_length]};
assign pixels_7_21 = {data_out[274*word_length-1 -: word_length]};
assign pixels_7_22 = {data_out[275*word_length-1 -: word_length]};
assign pixels_7_23 = {data_out[276*word_length-1 -: word_length]};
assign pixels_7_24 = {data_out[277*word_length-1 -: word_length]};
assign pixels_7_25 = {data_out[278*word_length-1 -: word_length]};
assign pixels_7_26 = {data_out[279*word_length-1 -: word_length]};
assign pixels_7_27 = {data_out[280*word_length-1 -: word_length]};
assign pixels_7_28 = {data_out[281*word_length-1 -: word_length]};
assign pixels_7_29 = {data_out[282*word_length-1 -: word_length]};
assign pixels_7_30 = {data_out[283*word_length-1 -: word_length]};
assign pixels_7_31 = {data_out[284*word_length-1 -: word_length]};
assign pixels_7_32 = {data_out[285*word_length-1 -: word_length]};
assign pixels_7_33 = {data_out[286*word_length-1 -: word_length]};
assign pixels_7_34 = {data_out[287*word_length-1 -: word_length]};
assign pixels_7_35 = {data_out[288*word_length-1 -: word_length]};
assign pixels_8_0 = {data_out[289*word_length-1 -: word_length]};
assign pixels_8_1 = {data_out[290*word_length-1 -: word_length]};
assign pixels_8_2 = {data_out[291*word_length-1 -: word_length]};
assign pixels_8_3 = {data_out[292*word_length-1 -: word_length]};
assign pixels_8_4 = {data_out[293*word_length-1 -: word_length]};
assign pixels_8_5 = {data_out[294*word_length-1 -: word_length]};
assign pixels_8_6 = {data_out[295*word_length-1 -: word_length]};
assign pixels_8_7 = {data_out[296*word_length-1 -: word_length]};
assign pixels_8_8 = {data_out[297*word_length-1 -: word_length]};
assign pixels_8_9 = {data_out[298*word_length-1 -: word_length]};
assign pixels_8_10 = {data_out[299*word_length-1 -: word_length]};
assign pixels_8_11 = {data_out[300*word_length-1 -: word_length]};
assign pixels_8_12 = {data_out[301*word_length-1 -: word_length]};
assign pixels_8_13 = {data_out[302*word_length-1 -: word_length]};
assign pixels_8_14 = {data_out[303*word_length-1 -: word_length]};
assign pixels_8_15 = {data_out[304*word_length-1 -: word_length]};
assign pixels_8_16 = {data_out[305*word_length-1 -: word_length]};
assign pixels_8_17 = {data_out[306*word_length-1 -: word_length]};
assign pixels_8_18 = {data_out[307*word_length-1 -: word_length]};
assign pixels_8_19 = {data_out[308*word_length-1 -: word_length]};
assign pixels_8_20 = {data_out[309*word_length-1 -: word_length]};
assign pixels_8_21 = {data_out[310*word_length-1 -: word_length]};
assign pixels_8_22 = {data_out[311*word_length-1 -: word_length]};
assign pixels_8_23 = {data_out[312*word_length-1 -: word_length]};
assign pixels_8_24 = {data_out[313*word_length-1 -: word_length]};
assign pixels_8_25 = {data_out[314*word_length-1 -: word_length]};
assign pixels_8_26 = {data_out[315*word_length-1 -: word_length]};
assign pixels_8_27 = {data_out[316*word_length-1 -: word_length]};
assign pixels_8_28 = {data_out[317*word_length-1 -: word_length]};
assign pixels_8_29 = {data_out[318*word_length-1 -: word_length]};
assign pixels_8_30 = {data_out[319*word_length-1 -: word_length]};
assign pixels_8_31 = {data_out[320*word_length-1 -: word_length]};
assign pixels_8_32 = {data_out[321*word_length-1 -: word_length]};
assign pixels_8_33 = {data_out[322*word_length-1 -: word_length]};
assign pixels_8_34 = {data_out[323*word_length-1 -: word_length]};
assign pixels_8_35 = {data_out[324*word_length-1 -: word_length]};
assign pixels_9_0 = {data_out[325*word_length-1 -: word_length]};
assign pixels_9_1 = {data_out[326*word_length-1 -: word_length]};
assign pixels_9_2 = {data_out[327*word_length-1 -: word_length]};
assign pixels_9_3 = {data_out[328*word_length-1 -: word_length]};
assign pixels_9_4 = {data_out[329*word_length-1 -: word_length]};
assign pixels_9_5 = {data_out[330*word_length-1 -: word_length]};
assign pixels_9_6 = {data_out[331*word_length-1 -: word_length]};
assign pixels_9_7 = {data_out[332*word_length-1 -: word_length]};
assign pixels_9_8 = {data_out[333*word_length-1 -: word_length]};
assign pixels_9_9 = {data_out[334*word_length-1 -: word_length]};
assign pixels_9_10 = {data_out[335*word_length-1 -: word_length]};
assign pixels_9_11 = {data_out[336*word_length-1 -: word_length]};
assign pixels_9_12 = {data_out[337*word_length-1 -: word_length]};
assign pixels_9_13 = {data_out[338*word_length-1 -: word_length]};
assign pixels_9_14 = {data_out[339*word_length-1 -: word_length]};
assign pixels_9_15 = {data_out[340*word_length-1 -: word_length]};
assign pixels_9_16 = {data_out[341*word_length-1 -: word_length]};
assign pixels_9_17 = {data_out[342*word_length-1 -: word_length]};
assign pixels_9_18 = {data_out[343*word_length-1 -: word_length]};
assign pixels_9_19 = {data_out[344*word_length-1 -: word_length]};
assign pixels_9_20 = {data_out[345*word_length-1 -: word_length]};
assign pixels_9_21 = {data_out[346*word_length-1 -: word_length]};
assign pixels_9_22 = {data_out[347*word_length-1 -: word_length]};
assign pixels_9_23 = {data_out[348*word_length-1 -: word_length]};
assign pixels_9_24 = {data_out[349*word_length-1 -: word_length]};
assign pixels_9_25 = {data_out[350*word_length-1 -: word_length]};
assign pixels_9_26 = {data_out[351*word_length-1 -: word_length]};
assign pixels_9_27 = {data_out[352*word_length-1 -: word_length]};
assign pixels_9_28 = {data_out[353*word_length-1 -: word_length]};
assign pixels_9_29 = {data_out[354*word_length-1 -: word_length]};
assign pixels_9_30 = {data_out[355*word_length-1 -: word_length]};
assign pixels_9_31 = {data_out[356*word_length-1 -: word_length]};
assign pixels_9_32 = {data_out[357*word_length-1 -: word_length]};
assign pixels_9_33 = {data_out[358*word_length-1 -: word_length]};
assign pixels_9_34 = {data_out[359*word_length-1 -: word_length]};
assign pixels_9_35 = {data_out[360*word_length-1 -: word_length]};
assign pixels_10_0 = {data_out[361*word_length-1 -: word_length]};
assign pixels_10_1 = {data_out[362*word_length-1 -: word_length]};
assign pixels_10_2 = {data_out[363*word_length-1 -: word_length]};
assign pixels_10_3 = {data_out[364*word_length-1 -: word_length]};
assign pixels_10_4 = {data_out[365*word_length-1 -: word_length]};
assign pixels_10_5 = {data_out[366*word_length-1 -: word_length]};
assign pixels_10_6 = {data_out[367*word_length-1 -: word_length]};
assign pixels_10_7 = {data_out[368*word_length-1 -: word_length]};
assign pixels_10_8 = {data_out[369*word_length-1 -: word_length]};
assign pixels_10_9 = {data_out[370*word_length-1 -: word_length]};
assign pixels_10_10 = {data_out[371*word_length-1 -: word_length]};
assign pixels_10_11 = {data_out[372*word_length-1 -: word_length]};
assign pixels_10_12 = {data_out[373*word_length-1 -: word_length]};
assign pixels_10_13 = {data_out[374*word_length-1 -: word_length]};
assign pixels_10_14 = {data_out[375*word_length-1 -: word_length]};
assign pixels_10_15 = {data_out[376*word_length-1 -: word_length]};
assign pixels_10_16 = {data_out[377*word_length-1 -: word_length]};
assign pixels_10_17 = {data_out[378*word_length-1 -: word_length]};
assign pixels_10_18 = {data_out[379*word_length-1 -: word_length]};
assign pixels_10_19 = {data_out[380*word_length-1 -: word_length]};
assign pixels_10_20 = {data_out[381*word_length-1 -: word_length]};
assign pixels_10_21 = {data_out[382*word_length-1 -: word_length]};
assign pixels_10_22 = {data_out[383*word_length-1 -: word_length]};
assign pixels_10_23 = {data_out[384*word_length-1 -: word_length]};
assign pixels_10_24 = {data_out[385*word_length-1 -: word_length]};
assign pixels_10_25 = {data_out[386*word_length-1 -: word_length]};
assign pixels_10_26 = {data_out[387*word_length-1 -: word_length]};
assign pixels_10_27 = {data_out[388*word_length-1 -: word_length]};
assign pixels_10_28 = {data_out[389*word_length-1 -: word_length]};
assign pixels_10_29 = {data_out[390*word_length-1 -: word_length]};
assign pixels_10_30 = {data_out[391*word_length-1 -: word_length]};
assign pixels_10_31 = {data_out[392*word_length-1 -: word_length]};
assign pixels_10_32 = {data_out[393*word_length-1 -: word_length]};
assign pixels_10_33 = {data_out[394*word_length-1 -: word_length]};
assign pixels_10_34 = {data_out[395*word_length-1 -: word_length]};
assign pixels_10_35 = {data_out[396*word_length-1 -: word_length]};
assign pixels_11_0 = {data_out[397*word_length-1 -: word_length]};
assign pixels_11_1 = {data_out[398*word_length-1 -: word_length]};
assign pixels_11_2 = {data_out[399*word_length-1 -: word_length]};
assign pixels_11_3 = {data_out[400*word_length-1 -: word_length]};
assign pixels_11_4 = {data_out[401*word_length-1 -: word_length]};
assign pixels_11_5 = {data_out[402*word_length-1 -: word_length]};
assign pixels_11_6 = {data_out[403*word_length-1 -: word_length]};
assign pixels_11_7 = {data_out[404*word_length-1 -: word_length]};
assign pixels_11_8 = {data_out[405*word_length-1 -: word_length]};
assign pixels_11_9 = {data_out[406*word_length-1 -: word_length]};
assign pixels_11_10 = {data_out[407*word_length-1 -: word_length]};
assign pixels_11_11 = {data_out[408*word_length-1 -: word_length]};
assign pixels_11_12 = {data_out[409*word_length-1 -: word_length]};
assign pixels_11_13 = {data_out[410*word_length-1 -: word_length]};
assign pixels_11_14 = {data_out[411*word_length-1 -: word_length]};
assign pixels_11_15 = {data_out[412*word_length-1 -: word_length]};
assign pixels_11_16 = {data_out[413*word_length-1 -: word_length]};
assign pixels_11_17 = {data_out[414*word_length-1 -: word_length]};
assign pixels_11_18 = {data_out[415*word_length-1 -: word_length]};
assign pixels_11_19 = {data_out[416*word_length-1 -: word_length]};
assign pixels_11_20 = {data_out[417*word_length-1 -: word_length]};
assign pixels_11_21 = {data_out[418*word_length-1 -: word_length]};
assign pixels_11_22 = {data_out[419*word_length-1 -: word_length]};
assign pixels_11_23 = {data_out[420*word_length-1 -: word_length]};
assign pixels_11_24 = {data_out[421*word_length-1 -: word_length]};
assign pixels_11_25 = {data_out[422*word_length-1 -: word_length]};
assign pixels_11_26 = {data_out[423*word_length-1 -: word_length]};
assign pixels_11_27 = {data_out[424*word_length-1 -: word_length]};
assign pixels_11_28 = {data_out[425*word_length-1 -: word_length]};
assign pixels_11_29 = {data_out[426*word_length-1 -: word_length]};
assign pixels_11_30 = {data_out[427*word_length-1 -: word_length]};
assign pixels_11_31 = {data_out[428*word_length-1 -: word_length]};
assign pixels_11_32 = {data_out[429*word_length-1 -: word_length]};
assign pixels_11_33 = {data_out[430*word_length-1 -: word_length]};
assign pixels_11_34 = {data_out[431*word_length-1 -: word_length]};
assign pixels_11_35 = {data_out[432*word_length-1 -: word_length]};
assign pixels_12_0 = {data_out[433*word_length-1 -: word_length]};
assign pixels_12_1 = {data_out[434*word_length-1 -: word_length]};
assign pixels_12_2 = {data_out[435*word_length-1 -: word_length]};
assign pixels_12_3 = {data_out[436*word_length-1 -: word_length]};
assign pixels_12_4 = {data_out[437*word_length-1 -: word_length]};
assign pixels_12_5 = {data_out[438*word_length-1 -: word_length]};
assign pixels_12_6 = {data_out[439*word_length-1 -: word_length]};
assign pixels_12_7 = {data_out[440*word_length-1 -: word_length]};
assign pixels_12_8 = {data_out[441*word_length-1 -: word_length]};
assign pixels_12_9 = {data_out[442*word_length-1 -: word_length]};
assign pixels_12_10 = {data_out[443*word_length-1 -: word_length]};
assign pixels_12_11 = {data_out[444*word_length-1 -: word_length]};
assign pixels_12_12 = {data_out[445*word_length-1 -: word_length]};
assign pixels_12_13 = {data_out[446*word_length-1 -: word_length]};
assign pixels_12_14 = {data_out[447*word_length-1 -: word_length]};
assign pixels_12_15 = {data_out[448*word_length-1 -: word_length]};
assign pixels_12_16 = {data_out[449*word_length-1 -: word_length]};
assign pixels_12_17 = {data_out[450*word_length-1 -: word_length]};
assign pixels_12_18 = {data_out[451*word_length-1 -: word_length]};
assign pixels_12_19 = {data_out[452*word_length-1 -: word_length]};
assign pixels_12_20 = {data_out[453*word_length-1 -: word_length]};
assign pixels_12_21 = {data_out[454*word_length-1 -: word_length]};
assign pixels_12_22 = {data_out[455*word_length-1 -: word_length]};
assign pixels_12_23 = {data_out[456*word_length-1 -: word_length]};
assign pixels_12_24 = {data_out[457*word_length-1 -: word_length]};
assign pixels_12_25 = {data_out[458*word_length-1 -: word_length]};
assign pixels_12_26 = {data_out[459*word_length-1 -: word_length]};
assign pixels_12_27 = {data_out[460*word_length-1 -: word_length]};
assign pixels_12_28 = {data_out[461*word_length-1 -: word_length]};
assign pixels_12_29 = {data_out[462*word_length-1 -: word_length]};
assign pixels_12_30 = {data_out[463*word_length-1 -: word_length]};
assign pixels_12_31 = {data_out[464*word_length-1 -: word_length]};
assign pixels_12_32 = {data_out[465*word_length-1 -: word_length]};
assign pixels_12_33 = {data_out[466*word_length-1 -: word_length]};
assign pixels_12_34 = {data_out[467*word_length-1 -: word_length]};
assign pixels_12_35 = {data_out[468*word_length-1 -: word_length]};
assign pixels_13_0 = {data_out[469*word_length-1 -: word_length]};
assign pixels_13_1 = {data_out[470*word_length-1 -: word_length]};
assign pixels_13_2 = {data_out[471*word_length-1 -: word_length]};
assign pixels_13_3 = {data_out[472*word_length-1 -: word_length]};
assign pixels_13_4 = {data_out[473*word_length-1 -: word_length]};
assign pixels_13_5 = {data_out[474*word_length-1 -: word_length]};
assign pixels_13_6 = {data_out[475*word_length-1 -: word_length]};
assign pixels_13_7 = {data_out[476*word_length-1 -: word_length]};
assign pixels_13_8 = {data_out[477*word_length-1 -: word_length]};
assign pixels_13_9 = {data_out[478*word_length-1 -: word_length]};
assign pixels_13_10 = {data_out[479*word_length-1 -: word_length]};
assign pixels_13_11 = {data_out[480*word_length-1 -: word_length]};
assign pixels_13_12 = {data_out[481*word_length-1 -: word_length]};
assign pixels_13_13 = {data_out[482*word_length-1 -: word_length]};
assign pixels_13_14 = {data_out[483*word_length-1 -: word_length]};
assign pixels_13_15 = {data_out[484*word_length-1 -: word_length]};
assign pixels_13_16 = {data_out[485*word_length-1 -: word_length]};
assign pixels_13_17 = {data_out[486*word_length-1 -: word_length]};
assign pixels_13_18 = {data_out[487*word_length-1 -: word_length]};
assign pixels_13_19 = {data_out[488*word_length-1 -: word_length]};
assign pixels_13_20 = {data_out[489*word_length-1 -: word_length]};
assign pixels_13_21 = {data_out[490*word_length-1 -: word_length]};
assign pixels_13_22 = {data_out[491*word_length-1 -: word_length]};
assign pixels_13_23 = {data_out[492*word_length-1 -: word_length]};
assign pixels_13_24 = {data_out[493*word_length-1 -: word_length]};
assign pixels_13_25 = {data_out[494*word_length-1 -: word_length]};
assign pixels_13_26 = {data_out[495*word_length-1 -: word_length]};
assign pixels_13_27 = {data_out[496*word_length-1 -: word_length]};
assign pixels_13_28 = {data_out[497*word_length-1 -: word_length]};
assign pixels_13_29 = {data_out[498*word_length-1 -: word_length]};
assign pixels_13_30 = {data_out[499*word_length-1 -: word_length]};
assign pixels_13_31 = {data_out[500*word_length-1 -: word_length]};
assign pixels_13_32 = {data_out[501*word_length-1 -: word_length]};
assign pixels_13_33 = {data_out[502*word_length-1 -: word_length]};
assign pixels_13_34 = {data_out[503*word_length-1 -: word_length]};
assign pixels_13_35 = {data_out[504*word_length-1 -: word_length]};
assign pixels_14_0 = {data_out[505*word_length-1 -: word_length]};
assign pixels_14_1 = {data_out[506*word_length-1 -: word_length]};
assign pixels_14_2 = {data_out[507*word_length-1 -: word_length]};
assign pixels_14_3 = {data_out[508*word_length-1 -: word_length]};
assign pixels_14_4 = {data_out[509*word_length-1 -: word_length]};
assign pixels_14_5 = {data_out[510*word_length-1 -: word_length]};
assign pixels_14_6 = {data_out[511*word_length-1 -: word_length]};
assign pixels_14_7 = {data_out[512*word_length-1 -: word_length]};
assign pixels_14_8 = {data_out[513*word_length-1 -: word_length]};
assign pixels_14_9 = {data_out[514*word_length-1 -: word_length]};
assign pixels_14_10 = {data_out[515*word_length-1 -: word_length]};
assign pixels_14_11 = {data_out[516*word_length-1 -: word_length]};
assign pixels_14_12 = {data_out[517*word_length-1 -: word_length]};
assign pixels_14_13 = {data_out[518*word_length-1 -: word_length]};
assign pixels_14_14 = {data_out[519*word_length-1 -: word_length]};
assign pixels_14_15 = {data_out[520*word_length-1 -: word_length]};
assign pixels_14_16 = {data_out[521*word_length-1 -: word_length]};
assign pixels_14_17 = {data_out[522*word_length-1 -: word_length]};
assign pixels_14_18 = {data_out[523*word_length-1 -: word_length]};
assign pixels_14_19 = {data_out[524*word_length-1 -: word_length]};
assign pixels_14_20 = {data_out[525*word_length-1 -: word_length]};
assign pixels_14_21 = {data_out[526*word_length-1 -: word_length]};
assign pixels_14_22 = {data_out[527*word_length-1 -: word_length]};
assign pixels_14_23 = {data_out[528*word_length-1 -: word_length]};
assign pixels_14_24 = {data_out[529*word_length-1 -: word_length]};
assign pixels_14_25 = {data_out[530*word_length-1 -: word_length]};
assign pixels_14_26 = {data_out[531*word_length-1 -: word_length]};
assign pixels_14_27 = {data_out[532*word_length-1 -: word_length]};
assign pixels_14_28 = {data_out[533*word_length-1 -: word_length]};
assign pixels_14_29 = {data_out[534*word_length-1 -: word_length]};
assign pixels_14_30 = {data_out[535*word_length-1 -: word_length]};
assign pixels_14_31 = {data_out[536*word_length-1 -: word_length]};
assign pixels_14_32 = {data_out[537*word_length-1 -: word_length]};
assign pixels_14_33 = {data_out[538*word_length-1 -: word_length]};
assign pixels_14_34 = {data_out[539*word_length-1 -: word_length]};
assign pixels_14_35 = {data_out[540*word_length-1 -: word_length]};
assign pixels_15_0 = {data_out[541*word_length-1 -: word_length]};
assign pixels_15_1 = {data_out[542*word_length-1 -: word_length]};
assign pixels_15_2 = {data_out[543*word_length-1 -: word_length]};
assign pixels_15_3 = {data_out[544*word_length-1 -: word_length]};
assign pixels_15_4 = {data_out[545*word_length-1 -: word_length]};
assign pixels_15_5 = {data_out[546*word_length-1 -: word_length]};
assign pixels_15_6 = {data_out[547*word_length-1 -: word_length]};
assign pixels_15_7 = {data_out[548*word_length-1 -: word_length]};
assign pixels_15_8 = {data_out[549*word_length-1 -: word_length]};
assign pixels_15_9 = {data_out[550*word_length-1 -: word_length]};
assign pixels_15_10 = {data_out[551*word_length-1 -: word_length]};
assign pixels_15_11 = {data_out[552*word_length-1 -: word_length]};
assign pixels_15_12 = {data_out[553*word_length-1 -: word_length]};
assign pixels_15_13 = {data_out[554*word_length-1 -: word_length]};
assign pixels_15_14 = {data_out[555*word_length-1 -: word_length]};
assign pixels_15_15 = {data_out[556*word_length-1 -: word_length]};
assign pixels_15_16 = {data_out[557*word_length-1 -: word_length]};
assign pixels_15_17 = {data_out[558*word_length-1 -: word_length]};
assign pixels_15_18 = {data_out[559*word_length-1 -: word_length]};
assign pixels_15_19 = {data_out[560*word_length-1 -: word_length]};
assign pixels_15_20 = {data_out[561*word_length-1 -: word_length]};
assign pixels_15_21 = {data_out[562*word_length-1 -: word_length]};
assign pixels_15_22 = {data_out[563*word_length-1 -: word_length]};
assign pixels_15_23 = {data_out[564*word_length-1 -: word_length]};
assign pixels_15_24 = {data_out[565*word_length-1 -: word_length]};
assign pixels_15_25 = {data_out[566*word_length-1 -: word_length]};
assign pixels_15_26 = {data_out[567*word_length-1 -: word_length]};
assign pixels_15_27 = {data_out[568*word_length-1 -: word_length]};
assign pixels_15_28 = {data_out[569*word_length-1 -: word_length]};
assign pixels_15_29 = {data_out[570*word_length-1 -: word_length]};
assign pixels_15_30 = {data_out[571*word_length-1 -: word_length]};
assign pixels_15_31 = {data_out[572*word_length-1 -: word_length]};
assign pixels_15_32 = {data_out[573*word_length-1 -: word_length]};
assign pixels_15_33 = {data_out[574*word_length-1 -: word_length]};
assign pixels_15_34 = {data_out[575*word_length-1 -: word_length]};
assign pixels_15_35 = {data_out[576*word_length-1 -: word_length]};
assign pixels_16_0 = {data_out[577*word_length-1 -: word_length]};
assign pixels_16_1 = {data_out[578*word_length-1 -: word_length]};
assign pixels_16_2 = {data_out[579*word_length-1 -: word_length]};
assign pixels_16_3 = {data_out[580*word_length-1 -: word_length]};
assign pixels_16_4 = {data_out[581*word_length-1 -: word_length]};
assign pixels_16_5 = {data_out[582*word_length-1 -: word_length]};
assign pixels_16_6 = {data_out[583*word_length-1 -: word_length]};
assign pixels_16_7 = {data_out[584*word_length-1 -: word_length]};
assign pixels_16_8 = {data_out[585*word_length-1 -: word_length]};
assign pixels_16_9 = {data_out[586*word_length-1 -: word_length]};
assign pixels_16_10 = {data_out[587*word_length-1 -: word_length]};
assign pixels_16_11 = {data_out[588*word_length-1 -: word_length]};
assign pixels_16_12 = {data_out[589*word_length-1 -: word_length]};
assign pixels_16_13 = {data_out[590*word_length-1 -: word_length]};
assign pixels_16_14 = {data_out[591*word_length-1 -: word_length]};
assign pixels_16_15 = {data_out[592*word_length-1 -: word_length]};
assign pixels_16_16 = {data_out[593*word_length-1 -: word_length]};
assign pixels_16_17 = {data_out[594*word_length-1 -: word_length]};
assign pixels_16_18 = {data_out[595*word_length-1 -: word_length]};
assign pixels_16_19 = {data_out[596*word_length-1 -: word_length]};
assign pixels_16_20 = {data_out[597*word_length-1 -: word_length]};
assign pixels_16_21 = {data_out[598*word_length-1 -: word_length]};
assign pixels_16_22 = {data_out[599*word_length-1 -: word_length]};
assign pixels_16_23 = {data_out[600*word_length-1 -: word_length]};
assign pixels_16_24 = {data_out[601*word_length-1 -: word_length]};
assign pixels_16_25 = {data_out[602*word_length-1 -: word_length]};
assign pixels_16_26 = {data_out[603*word_length-1 -: word_length]};
assign pixels_16_27 = {data_out[604*word_length-1 -: word_length]};
assign pixels_16_28 = {data_out[605*word_length-1 -: word_length]};
assign pixels_16_29 = {data_out[606*word_length-1 -: word_length]};
assign pixels_16_30 = {data_out[607*word_length-1 -: word_length]};
assign pixels_16_31 = {data_out[608*word_length-1 -: word_length]};
assign pixels_16_32 = {data_out[609*word_length-1 -: word_length]};
assign pixels_16_33 = {data_out[610*word_length-1 -: word_length]};
assign pixels_16_34 = {data_out[611*word_length-1 -: word_length]};
assign pixels_16_35 = {data_out[612*word_length-1 -: word_length]};
assign pixels_17_0 = {data_out[613*word_length-1 -: word_length]};
assign pixels_17_1 = {data_out[614*word_length-1 -: word_length]};
assign pixels_17_2 = {data_out[615*word_length-1 -: word_length]};
assign pixels_17_3 = {data_out[616*word_length-1 -: word_length]};
assign pixels_17_4 = {data_out[617*word_length-1 -: word_length]};
assign pixels_17_5 = {data_out[618*word_length-1 -: word_length]};
assign pixels_17_6 = {data_out[619*word_length-1 -: word_length]};
assign pixels_17_7 = {data_out[620*word_length-1 -: word_length]};
assign pixels_17_8 = {data_out[621*word_length-1 -: word_length]};
assign pixels_17_9 = {data_out[622*word_length-1 -: word_length]};
assign pixels_17_10 = {data_out[623*word_length-1 -: word_length]};
assign pixels_17_11 = {data_out[624*word_length-1 -: word_length]};
assign pixels_17_12 = {data_out[625*word_length-1 -: word_length]};
assign pixels_17_13 = {data_out[626*word_length-1 -: word_length]};
assign pixels_17_14 = {data_out[627*word_length-1 -: word_length]};
assign pixels_17_15 = {data_out[628*word_length-1 -: word_length]};
assign pixels_17_16 = {data_out[629*word_length-1 -: word_length]};
assign pixels_17_17 = {data_out[630*word_length-1 -: word_length]};
assign pixels_17_18 = {data_out[631*word_length-1 -: word_length]};
assign pixels_17_19 = {data_out[632*word_length-1 -: word_length]};
assign pixels_17_20 = {data_out[633*word_length-1 -: word_length]};
assign pixels_17_21 = {data_out[634*word_length-1 -: word_length]};
assign pixels_17_22 = {data_out[635*word_length-1 -: word_length]};
assign pixels_17_23 = {data_out[636*word_length-1 -: word_length]};
assign pixels_17_24 = {data_out[637*word_length-1 -: word_length]};
assign pixels_17_25 = {data_out[638*word_length-1 -: word_length]};
assign pixels_17_26 = {data_out[639*word_length-1 -: word_length]};
assign pixels_17_27 = {data_out[640*word_length-1 -: word_length]};
assign pixels_17_28 = {data_out[641*word_length-1 -: word_length]};
assign pixels_17_29 = {data_out[642*word_length-1 -: word_length]};
assign pixels_17_30 = {data_out[643*word_length-1 -: word_length]};
assign pixels_17_31 = {data_out[644*word_length-1 -: word_length]};
assign pixels_17_32 = {data_out[645*word_length-1 -: word_length]};
assign pixels_17_33 = {data_out[646*word_length-1 -: word_length]};
assign pixels_17_34 = {data_out[647*word_length-1 -: word_length]};
assign pixels_17_35 = {data_out[648*word_length-1 -: word_length]};
assign pixels_18_0 = {data_out[649*word_length-1 -: word_length]};
assign pixels_18_1 = {data_out[650*word_length-1 -: word_length]};
assign pixels_18_2 = {data_out[651*word_length-1 -: word_length]};
assign pixels_18_3 = {data_out[652*word_length-1 -: word_length]};
assign pixels_18_4 = {data_out[653*word_length-1 -: word_length]};
assign pixels_18_5 = {data_out[654*word_length-1 -: word_length]};
assign pixels_18_6 = {data_out[655*word_length-1 -: word_length]};
assign pixels_18_7 = {data_out[656*word_length-1 -: word_length]};
assign pixels_18_8 = {data_out[657*word_length-1 -: word_length]};
assign pixels_18_9 = {data_out[658*word_length-1 -: word_length]};
assign pixels_18_10 = {data_out[659*word_length-1 -: word_length]};
assign pixels_18_11 = {data_out[660*word_length-1 -: word_length]};
assign pixels_18_12 = {data_out[661*word_length-1 -: word_length]};
assign pixels_18_13 = {data_out[662*word_length-1 -: word_length]};
assign pixels_18_14 = {data_out[663*word_length-1 -: word_length]};
assign pixels_18_15 = {data_out[664*word_length-1 -: word_length]};
assign pixels_18_16 = {data_out[665*word_length-1 -: word_length]};
assign pixels_18_17 = {data_out[666*word_length-1 -: word_length]};
assign pixels_18_18 = {data_out[667*word_length-1 -: word_length]};
assign pixels_18_19 = {data_out[668*word_length-1 -: word_length]};
assign pixels_18_20 = {data_out[669*word_length-1 -: word_length]};
assign pixels_18_21 = {data_out[670*word_length-1 -: word_length]};
assign pixels_18_22 = {data_out[671*word_length-1 -: word_length]};
assign pixels_18_23 = {data_out[672*word_length-1 -: word_length]};
assign pixels_18_24 = {data_out[673*word_length-1 -: word_length]};
assign pixels_18_25 = {data_out[674*word_length-1 -: word_length]};
assign pixels_18_26 = {data_out[675*word_length-1 -: word_length]};
assign pixels_18_27 = {data_out[676*word_length-1 -: word_length]};
assign pixels_18_28 = {data_out[677*word_length-1 -: word_length]};
assign pixels_18_29 = {data_out[678*word_length-1 -: word_length]};
assign pixels_18_30 = {data_out[679*word_length-1 -: word_length]};
assign pixels_18_31 = {data_out[680*word_length-1 -: word_length]};
assign pixels_18_32 = {data_out[681*word_length-1 -: word_length]};
assign pixels_18_33 = {data_out[682*word_length-1 -: word_length]};
assign pixels_18_34 = {data_out[683*word_length-1 -: word_length]};
assign pixels_18_35 = {data_out[684*word_length-1 -: word_length]};
assign pixels_19_0 = {data_out[685*word_length-1 -: word_length]};
assign pixels_19_1 = {data_out[686*word_length-1 -: word_length]};
assign pixels_19_2 = {data_out[687*word_length-1 -: word_length]};
assign pixels_19_3 = {data_out[688*word_length-1 -: word_length]};
assign pixels_19_4 = {data_out[689*word_length-1 -: word_length]};
assign pixels_19_5 = {data_out[690*word_length-1 -: word_length]};
assign pixels_19_6 = {data_out[691*word_length-1 -: word_length]};
assign pixels_19_7 = {data_out[692*word_length-1 -: word_length]};
assign pixels_19_8 = {data_out[693*word_length-1 -: word_length]};
assign pixels_19_9 = {data_out[694*word_length-1 -: word_length]};
assign pixels_19_10 = {data_out[695*word_length-1 -: word_length]};
assign pixels_19_11 = {data_out[696*word_length-1 -: word_length]};
assign pixels_19_12 = {data_out[697*word_length-1 -: word_length]};
assign pixels_19_13 = {data_out[698*word_length-1 -: word_length]};
assign pixels_19_14 = {data_out[699*word_length-1 -: word_length]};
assign pixels_19_15 = {data_out[700*word_length-1 -: word_length]};
assign pixels_19_16 = {data_out[701*word_length-1 -: word_length]};
assign pixels_19_17 = {data_out[702*word_length-1 -: word_length]};
assign pixels_19_18 = {data_out[703*word_length-1 -: word_length]};
assign pixels_19_19 = {data_out[704*word_length-1 -: word_length]};
assign pixels_19_20 = {data_out[705*word_length-1 -: word_length]};
assign pixels_19_21 = {data_out[706*word_length-1 -: word_length]};
assign pixels_19_22 = {data_out[707*word_length-1 -: word_length]};
assign pixels_19_23 = {data_out[708*word_length-1 -: word_length]};
assign pixels_19_24 = {data_out[709*word_length-1 -: word_length]};
assign pixels_19_25 = {data_out[710*word_length-1 -: word_length]};
assign pixels_19_26 = {data_out[711*word_length-1 -: word_length]};
assign pixels_19_27 = {data_out[712*word_length-1 -: word_length]};
assign pixels_19_28 = {data_out[713*word_length-1 -: word_length]};
assign pixels_19_29 = {data_out[714*word_length-1 -: word_length]};
assign pixels_19_30 = {data_out[715*word_length-1 -: word_length]};
assign pixels_19_31 = {data_out[716*word_length-1 -: word_length]};
assign pixels_19_32 = {data_out[717*word_length-1 -: word_length]};
assign pixels_19_33 = {data_out[718*word_length-1 -: word_length]};
assign pixels_19_34 = {data_out[719*word_length-1 -: word_length]};
assign pixels_19_35 = {data_out[720*word_length-1 -: word_length]};
assign pixels_20_0 = {data_out[721*word_length-1 -: word_length]};
assign pixels_20_1 = {data_out[722*word_length-1 -: word_length]};
assign pixels_20_2 = {data_out[723*word_length-1 -: word_length]};
assign pixels_20_3 = {data_out[724*word_length-1 -: word_length]};
assign pixels_20_4 = {data_out[725*word_length-1 -: word_length]};
assign pixels_20_5 = {data_out[726*word_length-1 -: word_length]};
assign pixels_20_6 = {data_out[727*word_length-1 -: word_length]};
assign pixels_20_7 = {data_out[728*word_length-1 -: word_length]};
assign pixels_20_8 = {data_out[729*word_length-1 -: word_length]};
assign pixels_20_9 = {data_out[730*word_length-1 -: word_length]};
assign pixels_20_10 = {data_out[731*word_length-1 -: word_length]};
assign pixels_20_11 = {data_out[732*word_length-1 -: word_length]};
assign pixels_20_12 = {data_out[733*word_length-1 -: word_length]};
assign pixels_20_13 = {data_out[734*word_length-1 -: word_length]};
assign pixels_20_14 = {data_out[735*word_length-1 -: word_length]};
assign pixels_20_15 = {data_out[736*word_length-1 -: word_length]};
assign pixels_20_16 = {data_out[737*word_length-1 -: word_length]};
assign pixels_20_17 = {data_out[738*word_length-1 -: word_length]};
assign pixels_20_18 = {data_out[739*word_length-1 -: word_length]};
assign pixels_20_19 = {data_out[740*word_length-1 -: word_length]};
assign pixels_20_20 = {data_out[741*word_length-1 -: word_length]};
assign pixels_20_21 = {data_out[742*word_length-1 -: word_length]};
assign pixels_20_22 = {data_out[743*word_length-1 -: word_length]};
assign pixels_20_23 = {data_out[744*word_length-1 -: word_length]};
assign pixels_20_24 = {data_out[745*word_length-1 -: word_length]};
assign pixels_20_25 = {data_out[746*word_length-1 -: word_length]};
assign pixels_20_26 = {data_out[747*word_length-1 -: word_length]};
assign pixels_20_27 = {data_out[748*word_length-1 -: word_length]};
assign pixels_20_28 = {data_out[749*word_length-1 -: word_length]};
assign pixels_20_29 = {data_out[750*word_length-1 -: word_length]};
assign pixels_20_30 = {data_out[751*word_length-1 -: word_length]};
assign pixels_20_31 = {data_out[752*word_length-1 -: word_length]};
assign pixels_20_32 = {data_out[753*word_length-1 -: word_length]};
assign pixels_20_33 = {data_out[754*word_length-1 -: word_length]};
assign pixels_20_34 = {data_out[755*word_length-1 -: word_length]};
assign pixels_20_35 = {data_out[756*word_length-1 -: word_length]};
assign pixels_21_0 = {data_out[757*word_length-1 -: word_length]};
assign pixels_21_1 = {data_out[758*word_length-1 -: word_length]};
assign pixels_21_2 = {data_out[759*word_length-1 -: word_length]};
assign pixels_21_3 = {data_out[760*word_length-1 -: word_length]};
assign pixels_21_4 = {data_out[761*word_length-1 -: word_length]};
assign pixels_21_5 = {data_out[762*word_length-1 -: word_length]};
assign pixels_21_6 = {data_out[763*word_length-1 -: word_length]};
assign pixels_21_7 = {data_out[764*word_length-1 -: word_length]};
assign pixels_21_8 = {data_out[765*word_length-1 -: word_length]};
assign pixels_21_9 = {data_out[766*word_length-1 -: word_length]};
assign pixels_21_10 = {data_out[767*word_length-1 -: word_length]};
assign pixels_21_11 = {data_out[768*word_length-1 -: word_length]};
assign pixels_21_12 = {data_out[769*word_length-1 -: word_length]};
assign pixels_21_13 = {data_out[770*word_length-1 -: word_length]};
assign pixels_21_14 = {data_out[771*word_length-1 -: word_length]};
assign pixels_21_15 = {data_out[772*word_length-1 -: word_length]};
assign pixels_21_16 = {data_out[773*word_length-1 -: word_length]};
assign pixels_21_17 = {data_out[774*word_length-1 -: word_length]};
assign pixels_21_18 = {data_out[775*word_length-1 -: word_length]};
assign pixels_21_19 = {data_out[776*word_length-1 -: word_length]};
assign pixels_21_20 = {data_out[777*word_length-1 -: word_length]};
assign pixels_21_21 = {data_out[778*word_length-1 -: word_length]};
assign pixels_21_22 = {data_out[779*word_length-1 -: word_length]};
assign pixels_21_23 = {data_out[780*word_length-1 -: word_length]};
assign pixels_21_24 = {data_out[781*word_length-1 -: word_length]};
assign pixels_21_25 = {data_out[782*word_length-1 -: word_length]};
assign pixels_21_26 = {data_out[783*word_length-1 -: word_length]};
assign pixels_21_27 = {data_out[784*word_length-1 -: word_length]};
assign pixels_21_28 = {data_out[785*word_length-1 -: word_length]};
assign pixels_21_29 = {data_out[786*word_length-1 -: word_length]};
assign pixels_21_30 = {data_out[787*word_length-1 -: word_length]};
assign pixels_21_31 = {data_out[788*word_length-1 -: word_length]};
assign pixels_21_32 = {data_out[789*word_length-1 -: word_length]};
assign pixels_21_33 = {data_out[790*word_length-1 -: word_length]};
assign pixels_21_34 = {data_out[791*word_length-1 -: word_length]};
assign pixels_21_35 = {data_out[792*word_length-1 -: word_length]};
assign pixels_22_0 = {data_out[793*word_length-1 -: word_length]};
assign pixels_22_1 = {data_out[794*word_length-1 -: word_length]};
assign pixels_22_2 = {data_out[795*word_length-1 -: word_length]};
assign pixels_22_3 = {data_out[796*word_length-1 -: word_length]};
assign pixels_22_4 = {data_out[797*word_length-1 -: word_length]};
assign pixels_22_5 = {data_out[798*word_length-1 -: word_length]};
assign pixels_22_6 = {data_out[799*word_length-1 -: word_length]};
assign pixels_22_7 = {data_out[800*word_length-1 -: word_length]};
assign pixels_22_8 = {data_out[801*word_length-1 -: word_length]};
assign pixels_22_9 = {data_out[802*word_length-1 -: word_length]};
assign pixels_22_10 = {data_out[803*word_length-1 -: word_length]};
assign pixels_22_11 = {data_out[804*word_length-1 -: word_length]};
assign pixels_22_12 = {data_out[805*word_length-1 -: word_length]};
assign pixels_22_13 = {data_out[806*word_length-1 -: word_length]};
assign pixels_22_14 = {data_out[807*word_length-1 -: word_length]};
assign pixels_22_15 = {data_out[808*word_length-1 -: word_length]};
assign pixels_22_16 = {data_out[809*word_length-1 -: word_length]};
assign pixels_22_17 = {data_out[810*word_length-1 -: word_length]};
assign pixels_22_18 = {data_out[811*word_length-1 -: word_length]};
assign pixels_22_19 = {data_out[812*word_length-1 -: word_length]};
assign pixels_22_20 = {data_out[813*word_length-1 -: word_length]};
assign pixels_22_21 = {data_out[814*word_length-1 -: word_length]};
assign pixels_22_22 = {data_out[815*word_length-1 -: word_length]};
assign pixels_22_23 = {data_out[816*word_length-1 -: word_length]};
assign pixels_22_24 = {data_out[817*word_length-1 -: word_length]};
assign pixels_22_25 = {data_out[818*word_length-1 -: word_length]};
assign pixels_22_26 = {data_out[819*word_length-1 -: word_length]};
assign pixels_22_27 = {data_out[820*word_length-1 -: word_length]};
assign pixels_22_28 = {data_out[821*word_length-1 -: word_length]};
assign pixels_22_29 = {data_out[822*word_length-1 -: word_length]};
assign pixels_22_30 = {data_out[823*word_length-1 -: word_length]};
assign pixels_22_31 = {data_out[824*word_length-1 -: word_length]};
assign pixels_22_32 = {data_out[825*word_length-1 -: word_length]};
assign pixels_22_33 = {data_out[826*word_length-1 -: word_length]};
assign pixels_22_34 = {data_out[827*word_length-1 -: word_length]};
assign pixels_22_35 = {data_out[828*word_length-1 -: word_length]};
assign pixels_23_0 = {data_out[829*word_length-1 -: word_length]};
assign pixels_23_1 = {data_out[830*word_length-1 -: word_length]};
assign pixels_23_2 = {data_out[831*word_length-1 -: word_length]};
assign pixels_23_3 = {data_out[832*word_length-1 -: word_length]};
assign pixels_23_4 = {data_out[833*word_length-1 -: word_length]};
assign pixels_23_5 = {data_out[834*word_length-1 -: word_length]};
assign pixels_23_6 = {data_out[835*word_length-1 -: word_length]};
assign pixels_23_7 = {data_out[836*word_length-1 -: word_length]};
assign pixels_23_8 = {data_out[837*word_length-1 -: word_length]};
assign pixels_23_9 = {data_out[838*word_length-1 -: word_length]};
assign pixels_23_10 = {data_out[839*word_length-1 -: word_length]};
assign pixels_23_11 = {data_out[840*word_length-1 -: word_length]};
assign pixels_23_12 = {data_out[841*word_length-1 -: word_length]};
assign pixels_23_13 = {data_out[842*word_length-1 -: word_length]};
assign pixels_23_14 = {data_out[843*word_length-1 -: word_length]};
assign pixels_23_15 = {data_out[844*word_length-1 -: word_length]};
assign pixels_23_16 = {data_out[845*word_length-1 -: word_length]};
assign pixels_23_17 = {data_out[846*word_length-1 -: word_length]};
assign pixels_23_18 = {data_out[847*word_length-1 -: word_length]};
assign pixels_23_19 = {data_out[848*word_length-1 -: word_length]};
assign pixels_23_20 = {data_out[849*word_length-1 -: word_length]};
assign pixels_23_21 = {data_out[850*word_length-1 -: word_length]};
assign pixels_23_22 = {data_out[851*word_length-1 -: word_length]};
assign pixels_23_23 = {data_out[852*word_length-1 -: word_length]};
assign pixels_23_24 = {data_out[853*word_length-1 -: word_length]};
assign pixels_23_25 = {data_out[854*word_length-1 -: word_length]};
assign pixels_23_26 = {data_out[855*word_length-1 -: word_length]};
assign pixels_23_27 = {data_out[856*word_length-1 -: word_length]};
assign pixels_23_28 = {data_out[857*word_length-1 -: word_length]};
assign pixels_23_29 = {data_out[858*word_length-1 -: word_length]};
assign pixels_23_30 = {data_out[859*word_length-1 -: word_length]};
assign pixels_23_31 = {data_out[860*word_length-1 -: word_length]};
assign pixels_23_32 = {data_out[861*word_length-1 -: word_length]};
assign pixels_23_33 = {data_out[862*word_length-1 -: word_length]};
assign pixels_23_34 = {data_out[863*word_length-1 -: word_length]};
assign pixels_23_35 = {data_out[864*word_length-1 -: word_length]};
assign pixels_24_0 = {data_out[865*word_length-1 -: word_length]};
assign pixels_24_1 = {data_out[866*word_length-1 -: word_length]};
assign pixels_24_2 = {data_out[867*word_length-1 -: word_length]};
assign pixels_24_3 = {data_out[868*word_length-1 -: word_length]};
assign pixels_24_4 = {data_out[869*word_length-1 -: word_length]};
assign pixels_24_5 = {data_out[870*word_length-1 -: word_length]};
assign pixels_24_6 = {data_out[871*word_length-1 -: word_length]};
assign pixels_24_7 = {data_out[872*word_length-1 -: word_length]};
assign pixels_24_8 = {data_out[873*word_length-1 -: word_length]};
assign pixels_24_9 = {data_out[874*word_length-1 -: word_length]};
assign pixels_24_10 = {data_out[875*word_length-1 -: word_length]};
assign pixels_24_11 = {data_out[876*word_length-1 -: word_length]};
assign pixels_24_12 = {data_out[877*word_length-1 -: word_length]};
assign pixels_24_13 = {data_out[878*word_length-1 -: word_length]};
assign pixels_24_14 = {data_out[879*word_length-1 -: word_length]};
assign pixels_24_15 = {data_out[880*word_length-1 -: word_length]};
assign pixels_24_16 = {data_out[881*word_length-1 -: word_length]};
assign pixels_24_17 = {data_out[882*word_length-1 -: word_length]};
assign pixels_24_18 = {data_out[883*word_length-1 -: word_length]};
assign pixels_24_19 = {data_out[884*word_length-1 -: word_length]};
assign pixels_24_20 = {data_out[885*word_length-1 -: word_length]};
assign pixels_24_21 = {data_out[886*word_length-1 -: word_length]};
assign pixels_24_22 = {data_out[887*word_length-1 -: word_length]};
assign pixels_24_23 = {data_out[888*word_length-1 -: word_length]};
assign pixels_24_24 = {data_out[889*word_length-1 -: word_length]};
assign pixels_24_25 = {data_out[890*word_length-1 -: word_length]};
assign pixels_24_26 = {data_out[891*word_length-1 -: word_length]};
assign pixels_24_27 = {data_out[892*word_length-1 -: word_length]};
assign pixels_24_28 = {data_out[893*word_length-1 -: word_length]};
assign pixels_24_29 = {data_out[894*word_length-1 -: word_length]};
assign pixels_24_30 = {data_out[895*word_length-1 -: word_length]};
assign pixels_24_31 = {data_out[896*word_length-1 -: word_length]};
assign pixels_24_32 = {data_out[897*word_length-1 -: word_length]};
assign pixels_24_33 = {data_out[898*word_length-1 -: word_length]};
assign pixels_24_34 = {data_out[899*word_length-1 -: word_length]};
assign pixels_24_35 = {data_out[900*word_length-1 -: word_length]};
assign pixels_25_0 = {data_out[901*word_length-1 -: word_length]};
assign pixels_25_1 = {data_out[902*word_length-1 -: word_length]};
assign pixels_25_2 = {data_out[903*word_length-1 -: word_length]};
assign pixels_25_3 = {data_out[904*word_length-1 -: word_length]};
assign pixels_25_4 = {data_out[905*word_length-1 -: word_length]};
assign pixels_25_5 = {data_out[906*word_length-1 -: word_length]};
assign pixels_25_6 = {data_out[907*word_length-1 -: word_length]};
assign pixels_25_7 = {data_out[908*word_length-1 -: word_length]};
assign pixels_25_8 = {data_out[909*word_length-1 -: word_length]};
assign pixels_25_9 = {data_out[910*word_length-1 -: word_length]};
assign pixels_25_10 = {data_out[911*word_length-1 -: word_length]};
assign pixels_25_11 = {data_out[912*word_length-1 -: word_length]};
assign pixels_25_12 = {data_out[913*word_length-1 -: word_length]};
assign pixels_25_13 = {data_out[914*word_length-1 -: word_length]};
assign pixels_25_14 = {data_out[915*word_length-1 -: word_length]};
assign pixels_25_15 = {data_out[916*word_length-1 -: word_length]};
assign pixels_25_16 = {data_out[917*word_length-1 -: word_length]};
assign pixels_25_17 = {data_out[918*word_length-1 -: word_length]};
assign pixels_25_18 = {data_out[919*word_length-1 -: word_length]};
assign pixels_25_19 = {data_out[920*word_length-1 -: word_length]};
assign pixels_25_20 = {data_out[921*word_length-1 -: word_length]};
assign pixels_25_21 = {data_out[922*word_length-1 -: word_length]};
assign pixels_25_22 = {data_out[923*word_length-1 -: word_length]};
assign pixels_25_23 = {data_out[924*word_length-1 -: word_length]};
assign pixels_25_24 = {data_out[925*word_length-1 -: word_length]};
assign pixels_25_25 = {data_out[926*word_length-1 -: word_length]};
assign pixels_25_26 = {data_out[927*word_length-1 -: word_length]};
assign pixels_25_27 = {data_out[928*word_length-1 -: word_length]};
assign pixels_25_28 = {data_out[929*word_length-1 -: word_length]};
assign pixels_25_29 = {data_out[930*word_length-1 -: word_length]};
assign pixels_25_30 = {data_out[931*word_length-1 -: word_length]};
assign pixels_25_31 = {data_out[932*word_length-1 -: word_length]};
assign pixels_25_32 = {data_out[933*word_length-1 -: word_length]};
assign pixels_25_33 = {data_out[934*word_length-1 -: word_length]};
assign pixels_25_34 = {data_out[935*word_length-1 -: word_length]};
assign pixels_25_35 = {data_out[936*word_length-1 -: word_length]};
assign pixels_26_0 = {data_out[937*word_length-1 -: word_length]};
assign pixels_26_1 = {data_out[938*word_length-1 -: word_length]};
assign pixels_26_2 = {data_out[939*word_length-1 -: word_length]};
assign pixels_26_3 = {data_out[940*word_length-1 -: word_length]};
assign pixels_26_4 = {data_out[941*word_length-1 -: word_length]};
assign pixels_26_5 = {data_out[942*word_length-1 -: word_length]};
assign pixels_26_6 = {data_out[943*word_length-1 -: word_length]};
assign pixels_26_7 = {data_out[944*word_length-1 -: word_length]};
assign pixels_26_8 = {data_out[945*word_length-1 -: word_length]};
assign pixels_26_9 = {data_out[946*word_length-1 -: word_length]};
assign pixels_26_10 = {data_out[947*word_length-1 -: word_length]};
assign pixels_26_11 = {data_out[948*word_length-1 -: word_length]};
assign pixels_26_12 = {data_out[949*word_length-1 -: word_length]};
assign pixels_26_13 = {data_out[950*word_length-1 -: word_length]};
assign pixels_26_14 = {data_out[951*word_length-1 -: word_length]};
assign pixels_26_15 = {data_out[952*word_length-1 -: word_length]};
assign pixels_26_16 = {data_out[953*word_length-1 -: word_length]};
assign pixels_26_17 = {data_out[954*word_length-1 -: word_length]};
assign pixels_26_18 = {data_out[955*word_length-1 -: word_length]};
assign pixels_26_19 = {data_out[956*word_length-1 -: word_length]};
assign pixels_26_20 = {data_out[957*word_length-1 -: word_length]};
assign pixels_26_21 = {data_out[958*word_length-1 -: word_length]};
assign pixels_26_22 = {data_out[959*word_length-1 -: word_length]};
assign pixels_26_23 = {data_out[960*word_length-1 -: word_length]};
assign pixels_26_24 = {data_out[961*word_length-1 -: word_length]};
assign pixels_26_25 = {data_out[962*word_length-1 -: word_length]};
assign pixels_26_26 = {data_out[963*word_length-1 -: word_length]};
assign pixels_26_27 = {data_out[964*word_length-1 -: word_length]};
assign pixels_26_28 = {data_out[965*word_length-1 -: word_length]};
assign pixels_26_29 = {data_out[966*word_length-1 -: word_length]};
assign pixels_26_30 = {data_out[967*word_length-1 -: word_length]};
assign pixels_26_31 = {data_out[968*word_length-1 -: word_length]};
assign pixels_26_32 = {data_out[969*word_length-1 -: word_length]};
assign pixels_26_33 = {data_out[970*word_length-1 -: word_length]};
assign pixels_26_34 = {data_out[971*word_length-1 -: word_length]};
assign pixels_26_35 = {data_out[972*word_length-1 -: word_length]};
assign pixels_27_0 = {data_out[973*word_length-1 -: word_length]};
assign pixels_27_1 = {data_out[974*word_length-1 -: word_length]};
assign pixels_27_2 = {data_out[975*word_length-1 -: word_length]};
assign pixels_27_3 = {data_out[976*word_length-1 -: word_length]};
assign pixels_27_4 = {data_out[977*word_length-1 -: word_length]};
assign pixels_27_5 = {data_out[978*word_length-1 -: word_length]};
assign pixels_27_6 = {data_out[979*word_length-1 -: word_length]};
assign pixels_27_7 = {data_out[980*word_length-1 -: word_length]};
assign pixels_27_8 = {data_out[981*word_length-1 -: word_length]};
assign pixels_27_9 = {data_out[982*word_length-1 -: word_length]};
assign pixels_27_10 = {data_out[983*word_length-1 -: word_length]};
assign pixels_27_11 = {data_out[984*word_length-1 -: word_length]};
assign pixels_27_12 = {data_out[985*word_length-1 -: word_length]};
assign pixels_27_13 = {data_out[986*word_length-1 -: word_length]};
assign pixels_27_14 = {data_out[987*word_length-1 -: word_length]};
assign pixels_27_15 = {data_out[988*word_length-1 -: word_length]};
assign pixels_27_16 = {data_out[989*word_length-1 -: word_length]};
assign pixels_27_17 = {data_out[990*word_length-1 -: word_length]};
assign pixels_27_18 = {data_out[991*word_length-1 -: word_length]};
assign pixels_27_19 = {data_out[992*word_length-1 -: word_length]};
assign pixels_27_20 = {data_out[993*word_length-1 -: word_length]};
assign pixels_27_21 = {data_out[994*word_length-1 -: word_length]};
assign pixels_27_22 = {data_out[995*word_length-1 -: word_length]};
assign pixels_27_23 = {data_out[996*word_length-1 -: word_length]};
assign pixels_27_24 = {data_out[997*word_length-1 -: word_length]};
assign pixels_27_25 = {data_out[998*word_length-1 -: word_length]};
assign pixels_27_26 = {data_out[999*word_length-1 -: word_length]};
assign pixels_27_27 = {data_out[1000*word_length-1 -: word_length]};
assign pixels_27_28 = {data_out[1001*word_length-1 -: word_length]};
assign pixels_27_29 = {data_out[1002*word_length-1 -: word_length]};
assign pixels_27_30 = {data_out[1003*word_length-1 -: word_length]};
assign pixels_27_31 = {data_out[1004*word_length-1 -: word_length]};
assign pixels_27_32 = {data_out[1005*word_length-1 -: word_length]};
assign pixels_27_33 = {data_out[1006*word_length-1 -: word_length]};
assign pixels_27_34 = {data_out[1007*word_length-1 -: word_length]};
assign pixels_27_35 = {data_out[1008*word_length-1 -: word_length]};
assign pixels_28_0 = {data_out[1009*word_length-1 -: word_length]};
assign pixels_28_1 = {data_out[1010*word_length-1 -: word_length]};
assign pixels_28_2 = {data_out[1011*word_length-1 -: word_length]};
assign pixels_28_3 = {data_out[1012*word_length-1 -: word_length]};
assign pixels_28_4 = {data_out[1013*word_length-1 -: word_length]};
assign pixels_28_5 = {data_out[1014*word_length-1 -: word_length]};
assign pixels_28_6 = {data_out[1015*word_length-1 -: word_length]};
assign pixels_28_7 = {data_out[1016*word_length-1 -: word_length]};
assign pixels_28_8 = {data_out[1017*word_length-1 -: word_length]};
assign pixels_28_9 = {data_out[1018*word_length-1 -: word_length]};
assign pixels_28_10 = {data_out[1019*word_length-1 -: word_length]};
assign pixels_28_11 = {data_out[1020*word_length-1 -: word_length]};
assign pixels_28_12 = {data_out[1021*word_length-1 -: word_length]};
assign pixels_28_13 = {data_out[1022*word_length-1 -: word_length]};
assign pixels_28_14 = {data_out[1023*word_length-1 -: word_length]};
assign pixels_28_15 = {data_out[1024*word_length-1 -: word_length]};
assign pixels_28_16 = {data_out[1025*word_length-1 -: word_length]};
assign pixels_28_17 = {data_out[1026*word_length-1 -: word_length]};
assign pixels_28_18 = {data_out[1027*word_length-1 -: word_length]};
assign pixels_28_19 = {data_out[1028*word_length-1 -: word_length]};
assign pixels_28_20 = {data_out[1029*word_length-1 -: word_length]};
assign pixels_28_21 = {data_out[1030*word_length-1 -: word_length]};
assign pixels_28_22 = {data_out[1031*word_length-1 -: word_length]};
assign pixels_28_23 = {data_out[1032*word_length-1 -: word_length]};
assign pixels_28_24 = {data_out[1033*word_length-1 -: word_length]};
assign pixels_28_25 = {data_out[1034*word_length-1 -: word_length]};
assign pixels_28_26 = {data_out[1035*word_length-1 -: word_length]};
assign pixels_28_27 = {data_out[1036*word_length-1 -: word_length]};
assign pixels_28_28 = {data_out[1037*word_length-1 -: word_length]};
assign pixels_28_29 = {data_out[1038*word_length-1 -: word_length]};
assign pixels_28_30 = {data_out[1039*word_length-1 -: word_length]};
assign pixels_28_31 = {data_out[1040*word_length-1 -: word_length]};
assign pixels_28_32 = {data_out[1041*word_length-1 -: word_length]};
assign pixels_28_33 = {data_out[1042*word_length-1 -: word_length]};
assign pixels_28_34 = {data_out[1043*word_length-1 -: word_length]};
assign pixels_28_35 = {data_out[1044*word_length-1 -: word_length]};
assign pixels_29_0 = {data_out[1045*word_length-1 -: word_length]};
assign pixels_29_1 = {data_out[1046*word_length-1 -: word_length]};
assign pixels_29_2 = {data_out[1047*word_length-1 -: word_length]};
assign pixels_29_3 = {data_out[1048*word_length-1 -: word_length]};
assign pixels_29_4 = {data_out[1049*word_length-1 -: word_length]};
assign pixels_29_5 = {data_out[1050*word_length-1 -: word_length]};
assign pixels_29_6 = {data_out[1051*word_length-1 -: word_length]};
assign pixels_29_7 = {data_out[1052*word_length-1 -: word_length]};
assign pixels_29_8 = {data_out[1053*word_length-1 -: word_length]};
assign pixels_29_9 = {data_out[1054*word_length-1 -: word_length]};
assign pixels_29_10 = {data_out[1055*word_length-1 -: word_length]};
assign pixels_29_11 = {data_out[1056*word_length-1 -: word_length]};
assign pixels_29_12 = {data_out[1057*word_length-1 -: word_length]};
assign pixels_29_13 = {data_out[1058*word_length-1 -: word_length]};
assign pixels_29_14 = {data_out[1059*word_length-1 -: word_length]};
assign pixels_29_15 = {data_out[1060*word_length-1 -: word_length]};
assign pixels_29_16 = {data_out[1061*word_length-1 -: word_length]};
assign pixels_29_17 = {data_out[1062*word_length-1 -: word_length]};
assign pixels_29_18 = {data_out[1063*word_length-1 -: word_length]};
assign pixels_29_19 = {data_out[1064*word_length-1 -: word_length]};
assign pixels_29_20 = {data_out[1065*word_length-1 -: word_length]};
assign pixels_29_21 = {data_out[1066*word_length-1 -: word_length]};
assign pixels_29_22 = {data_out[1067*word_length-1 -: word_length]};
assign pixels_29_23 = {data_out[1068*word_length-1 -: word_length]};
assign pixels_29_24 = {data_out[1069*word_length-1 -: word_length]};
assign pixels_29_25 = {data_out[1070*word_length-1 -: word_length]};
assign pixels_29_26 = {data_out[1071*word_length-1 -: word_length]};
assign pixels_29_27 = {data_out[1072*word_length-1 -: word_length]};
assign pixels_29_28 = {data_out[1073*word_length-1 -: word_length]};
assign pixels_29_29 = {data_out[1074*word_length-1 -: word_length]};
assign pixels_29_30 = {data_out[1075*word_length-1 -: word_length]};
assign pixels_29_31 = {data_out[1076*word_length-1 -: word_length]};
assign pixels_29_32 = {data_out[1077*word_length-1 -: word_length]};
assign pixels_29_33 = {data_out[1078*word_length-1 -: word_length]};
assign pixels_29_34 = {data_out[1079*word_length-1 -: word_length]};
assign pixels_29_35 = {data_out[1080*word_length-1 -: word_length]};
assign pixels_30_0 = {data_out[1081*word_length-1 -: word_length]};
assign pixels_30_1 = {data_out[1082*word_length-1 -: word_length]};
assign pixels_30_2 = {data_out[1083*word_length-1 -: word_length]};
assign pixels_30_3 = {data_out[1084*word_length-1 -: word_length]};
assign pixels_30_4 = {data_out[1085*word_length-1 -: word_length]};
assign pixels_30_5 = {data_out[1086*word_length-1 -: word_length]};
assign pixels_30_6 = {data_out[1087*word_length-1 -: word_length]};
assign pixels_30_7 = {data_out[1088*word_length-1 -: word_length]};
assign pixels_30_8 = {data_out[1089*word_length-1 -: word_length]};
assign pixels_30_9 = {data_out[1090*word_length-1 -: word_length]};
assign pixels_30_10 = {data_out[1091*word_length-1 -: word_length]};
assign pixels_30_11 = {data_out[1092*word_length-1 -: word_length]};
assign pixels_30_12 = {data_out[1093*word_length-1 -: word_length]};
assign pixels_30_13 = {data_out[1094*word_length-1 -: word_length]};
assign pixels_30_14 = {data_out[1095*word_length-1 -: word_length]};
assign pixels_30_15 = {data_out[1096*word_length-1 -: word_length]};
assign pixels_30_16 = {data_out[1097*word_length-1 -: word_length]};
assign pixels_30_17 = {data_out[1098*word_length-1 -: word_length]};
assign pixels_30_18 = {data_out[1099*word_length-1 -: word_length]};
assign pixels_30_19 = {data_out[1100*word_length-1 -: word_length]};
assign pixels_30_20 = {data_out[1101*word_length-1 -: word_length]};
assign pixels_30_21 = {data_out[1102*word_length-1 -: word_length]};
assign pixels_30_22 = {data_out[1103*word_length-1 -: word_length]};
assign pixels_30_23 = {data_out[1104*word_length-1 -: word_length]};
assign pixels_30_24 = {data_out[1105*word_length-1 -: word_length]};
assign pixels_30_25 = {data_out[1106*word_length-1 -: word_length]};
assign pixels_30_26 = {data_out[1107*word_length-1 -: word_length]};
assign pixels_30_27 = {data_out[1108*word_length-1 -: word_length]};
assign pixels_30_28 = {data_out[1109*word_length-1 -: word_length]};
assign pixels_30_29 = {data_out[1110*word_length-1 -: word_length]};
assign pixels_30_30 = {data_out[1111*word_length-1 -: word_length]};
assign pixels_30_31 = {data_out[1112*word_length-1 -: word_length]};
assign pixels_30_32 = {data_out[1113*word_length-1 -: word_length]};
assign pixels_30_33 = {data_out[1114*word_length-1 -: word_length]};
assign pixels_30_34 = {data_out[1115*word_length-1 -: word_length]};
assign pixels_30_35 = {data_out[1116*word_length-1 -: word_length]};
assign pixels_31_0 = {data_out[1117*word_length-1 -: word_length]};
assign pixels_31_1 = {data_out[1118*word_length-1 -: word_length]};
assign pixels_31_2 = {data_out[1119*word_length-1 -: word_length]};
assign pixels_31_3 = {data_out[1120*word_length-1 -: word_length]};
assign pixels_31_4 = {data_out[1121*word_length-1 -: word_length]};
assign pixels_31_5 = {data_out[1122*word_length-1 -: word_length]};
assign pixels_31_6 = {data_out[1123*word_length-1 -: word_length]};
assign pixels_31_7 = {data_out[1124*word_length-1 -: word_length]};
assign pixels_31_8 = {data_out[1125*word_length-1 -: word_length]};
assign pixels_31_9 = {data_out[1126*word_length-1 -: word_length]};
assign pixels_31_10 = {data_out[1127*word_length-1 -: word_length]};
assign pixels_31_11 = {data_out[1128*word_length-1 -: word_length]};
assign pixels_31_12 = {data_out[1129*word_length-1 -: word_length]};
assign pixels_31_13 = {data_out[1130*word_length-1 -: word_length]};
assign pixels_31_14 = {data_out[1131*word_length-1 -: word_length]};
assign pixels_31_15 = {data_out[1132*word_length-1 -: word_length]};
assign pixels_31_16 = {data_out[1133*word_length-1 -: word_length]};
assign pixels_31_17 = {data_out[1134*word_length-1 -: word_length]};
assign pixels_31_18 = {data_out[1135*word_length-1 -: word_length]};
assign pixels_31_19 = {data_out[1136*word_length-1 -: word_length]};
assign pixels_31_20 = {data_out[1137*word_length-1 -: word_length]};
assign pixels_31_21 = {data_out[1138*word_length-1 -: word_length]};
assign pixels_31_22 = {data_out[1139*word_length-1 -: word_length]};
assign pixels_31_23 = {data_out[1140*word_length-1 -: word_length]};
assign pixels_31_24 = {data_out[1141*word_length-1 -: word_length]};
assign pixels_31_25 = {data_out[1142*word_length-1 -: word_length]};
assign pixels_31_26 = {data_out[1143*word_length-1 -: word_length]};
assign pixels_31_27 = {data_out[1144*word_length-1 -: word_length]};
assign pixels_31_28 = {data_out[1145*word_length-1 -: word_length]};
assign pixels_31_29 = {data_out[1146*word_length-1 -: word_length]};
assign pixels_31_30 = {data_out[1147*word_length-1 -: word_length]};
assign pixels_31_31 = {data_out[1148*word_length-1 -: word_length]};
assign pixels_31_32 = {data_out[1149*word_length-1 -: word_length]};
assign pixels_31_33 = {data_out[1150*word_length-1 -: word_length]};
assign pixels_31_34 = {data_out[1151*word_length-1 -: word_length]};
assign pixels_31_35 = {data_out[1152*word_length-1 -: word_length]};
assign pixels_32_0 = {data_out[1153*word_length-1 -: word_length]};
assign pixels_32_1 = {data_out[1154*word_length-1 -: word_length]};
assign pixels_32_2 = {data_out[1155*word_length-1 -: word_length]};
assign pixels_32_3 = {data_out[1156*word_length-1 -: word_length]};
assign pixels_32_4 = {data_out[1157*word_length-1 -: word_length]};
assign pixels_32_5 = {data_out[1158*word_length-1 -: word_length]};
assign pixels_32_6 = {data_out[1159*word_length-1 -: word_length]};
assign pixels_32_7 = {data_out[1160*word_length-1 -: word_length]};
assign pixels_32_8 = {data_out[1161*word_length-1 -: word_length]};
assign pixels_32_9 = {data_out[1162*word_length-1 -: word_length]};
assign pixels_32_10 = {data_out[1163*word_length-1 -: word_length]};
assign pixels_32_11 = {data_out[1164*word_length-1 -: word_length]};
assign pixels_32_12 = {data_out[1165*word_length-1 -: word_length]};
assign pixels_32_13 = {data_out[1166*word_length-1 -: word_length]};
assign pixels_32_14 = {data_out[1167*word_length-1 -: word_length]};
assign pixels_32_15 = {data_out[1168*word_length-1 -: word_length]};
assign pixels_32_16 = {data_out[1169*word_length-1 -: word_length]};
assign pixels_32_17 = {data_out[1170*word_length-1 -: word_length]};
assign pixels_32_18 = {data_out[1171*word_length-1 -: word_length]};
assign pixels_32_19 = {data_out[1172*word_length-1 -: word_length]};
assign pixels_32_20 = {data_out[1173*word_length-1 -: word_length]};
assign pixels_32_21 = {data_out[1174*word_length-1 -: word_length]};
assign pixels_32_22 = {data_out[1175*word_length-1 -: word_length]};
assign pixels_32_23 = {data_out[1176*word_length-1 -: word_length]};
assign pixels_32_24 = {data_out[1177*word_length-1 -: word_length]};
assign pixels_32_25 = {data_out[1178*word_length-1 -: word_length]};
assign pixels_32_26 = {data_out[1179*word_length-1 -: word_length]};
assign pixels_32_27 = {data_out[1180*word_length-1 -: word_length]};
assign pixels_32_28 = {data_out[1181*word_length-1 -: word_length]};
assign pixels_32_29 = {data_out[1182*word_length-1 -: word_length]};
assign pixels_32_30 = {data_out[1183*word_length-1 -: word_length]};
assign pixels_32_31 = {data_out[1184*word_length-1 -: word_length]};
assign pixels_32_32 = {data_out[1185*word_length-1 -: word_length]};
assign pixels_32_33 = {data_out[1186*word_length-1 -: word_length]};
assign pixels_32_34 = {data_out[1187*word_length-1 -: word_length]};
assign pixels_32_35 = {data_out[1188*word_length-1 -: word_length]};
assign pixels_33_0 = {data_out[1189*word_length-1 -: word_length]};
assign pixels_33_1 = {data_out[1190*word_length-1 -: word_length]};
assign pixels_33_2 = {data_out[1191*word_length-1 -: word_length]};
assign pixels_33_3 = {data_out[1192*word_length-1 -: word_length]};
assign pixels_33_4 = {data_out[1193*word_length-1 -: word_length]};
assign pixels_33_5 = {data_out[1194*word_length-1 -: word_length]};
assign pixels_33_6 = {data_out[1195*word_length-1 -: word_length]};
assign pixels_33_7 = {data_out[1196*word_length-1 -: word_length]};
assign pixels_33_8 = {data_out[1197*word_length-1 -: word_length]};
assign pixels_33_9 = {data_out[1198*word_length-1 -: word_length]};
assign pixels_33_10 = {data_out[1199*word_length-1 -: word_length]};
assign pixels_33_11 = {data_out[1200*word_length-1 -: word_length]};
assign pixels_33_12 = {data_out[1201*word_length-1 -: word_length]};
assign pixels_33_13 = {data_out[1202*word_length-1 -: word_length]};
assign pixels_33_14 = {data_out[1203*word_length-1 -: word_length]};
assign pixels_33_15 = {data_out[1204*word_length-1 -: word_length]};
assign pixels_33_16 = {data_out[1205*word_length-1 -: word_length]};
assign pixels_33_17 = {data_out[1206*word_length-1 -: word_length]};
assign pixels_33_18 = {data_out[1207*word_length-1 -: word_length]};
assign pixels_33_19 = {data_out[1208*word_length-1 -: word_length]};
assign pixels_33_20 = {data_out[1209*word_length-1 -: word_length]};
assign pixels_33_21 = {data_out[1210*word_length-1 -: word_length]};
assign pixels_33_22 = {data_out[1211*word_length-1 -: word_length]};
assign pixels_33_23 = {data_out[1212*word_length-1 -: word_length]};
assign pixels_33_24 = {data_out[1213*word_length-1 -: word_length]};
assign pixels_33_25 = {data_out[1214*word_length-1 -: word_length]};
assign pixels_33_26 = {data_out[1215*word_length-1 -: word_length]};
assign pixels_33_27 = {data_out[1216*word_length-1 -: word_length]};
assign pixels_33_28 = {data_out[1217*word_length-1 -: word_length]};
assign pixels_33_29 = {data_out[1218*word_length-1 -: word_length]};
assign pixels_33_30 = {data_out[1219*word_length-1 -: word_length]};
assign pixels_33_31 = {data_out[1220*word_length-1 -: word_length]};
assign pixels_33_32 = {data_out[1221*word_length-1 -: word_length]};
assign pixels_33_33 = {data_out[1222*word_length-1 -: word_length]};
assign pixels_33_34 = {data_out[1223*word_length-1 -: word_length]};
assign pixels_33_35 = {data_out[1224*word_length-1 -: word_length]};
assign pixels_34_0 = {data_out[1225*word_length-1 -: word_length]};
assign pixels_34_1 = {data_out[1226*word_length-1 -: word_length]};
assign pixels_34_2 = {data_out[1227*word_length-1 -: word_length]};
assign pixels_34_3 = {data_out[1228*word_length-1 -: word_length]};
assign pixels_34_4 = {data_out[1229*word_length-1 -: word_length]};
assign pixels_34_5 = {data_out[1230*word_length-1 -: word_length]};
assign pixels_34_6 = {data_out[1231*word_length-1 -: word_length]};
assign pixels_34_7 = {data_out[1232*word_length-1 -: word_length]};
assign pixels_34_8 = {data_out[1233*word_length-1 -: word_length]};
assign pixels_34_9 = {data_out[1234*word_length-1 -: word_length]};
assign pixels_34_10 = {data_out[1235*word_length-1 -: word_length]};
assign pixels_34_11 = {data_out[1236*word_length-1 -: word_length]};
assign pixels_34_12 = {data_out[1237*word_length-1 -: word_length]};
assign pixels_34_13 = {data_out[1238*word_length-1 -: word_length]};
assign pixels_34_14 = {data_out[1239*word_length-1 -: word_length]};
assign pixels_34_15 = {data_out[1240*word_length-1 -: word_length]};
assign pixels_34_16 = {data_out[1241*word_length-1 -: word_length]};
assign pixels_34_17 = {data_out[1242*word_length-1 -: word_length]};
assign pixels_34_18 = {data_out[1243*word_length-1 -: word_length]};
assign pixels_34_19 = {data_out[1244*word_length-1 -: word_length]};
assign pixels_34_20 = {data_out[1245*word_length-1 -: word_length]};
assign pixels_34_21 = {data_out[1246*word_length-1 -: word_length]};
assign pixels_34_22 = {data_out[1247*word_length-1 -: word_length]};
assign pixels_34_23 = {data_out[1248*word_length-1 -: word_length]};
assign pixels_34_24 = {data_out[1249*word_length-1 -: word_length]};
assign pixels_34_25 = {data_out[1250*word_length-1 -: word_length]};
assign pixels_34_26 = {data_out[1251*word_length-1 -: word_length]};
assign pixels_34_27 = {data_out[1252*word_length-1 -: word_length]};
assign pixels_34_28 = {data_out[1253*word_length-1 -: word_length]};
assign pixels_34_29 = {data_out[1254*word_length-1 -: word_length]};
assign pixels_34_30 = {data_out[1255*word_length-1 -: word_length]};
assign pixels_34_31 = {data_out[1256*word_length-1 -: word_length]};
assign pixels_34_32 = {data_out[1257*word_length-1 -: word_length]};
assign pixels_34_33 = {data_out[1258*word_length-1 -: word_length]};
assign pixels_34_34 = {data_out[1259*word_length-1 -: word_length]};
assign pixels_34_35 = {data_out[1260*word_length-1 -: word_length]};
assign pixels_35_0 = {data_out[1261*word_length-1 -: word_length]};
assign pixels_35_1 = {data_out[1262*word_length-1 -: word_length]};
assign pixels_35_2 = {data_out[1263*word_length-1 -: word_length]};
assign pixels_35_3 = {data_out[1264*word_length-1 -: word_length]};
assign pixels_35_4 = {data_out[1265*word_length-1 -: word_length]};
assign pixels_35_5 = {data_out[1266*word_length-1 -: word_length]};
assign pixels_35_6 = {data_out[1267*word_length-1 -: word_length]};
assign pixels_35_7 = {data_out[1268*word_length-1 -: word_length]};
assign pixels_35_8 = {data_out[1269*word_length-1 -: word_length]};
assign pixels_35_9 = {data_out[1270*word_length-1 -: word_length]};
assign pixels_35_10 = {data_out[1271*word_length-1 -: word_length]};
assign pixels_35_11 = {data_out[1272*word_length-1 -: word_length]};
assign pixels_35_12 = {data_out[1273*word_length-1 -: word_length]};
assign pixels_35_13 = {data_out[1274*word_length-1 -: word_length]};
assign pixels_35_14 = {data_out[1275*word_length-1 -: word_length]};
assign pixels_35_15 = {data_out[1276*word_length-1 -: word_length]};
assign pixels_35_16 = {data_out[1277*word_length-1 -: word_length]};
assign pixels_35_17 = {data_out[1278*word_length-1 -: word_length]};
assign pixels_35_18 = {data_out[1279*word_length-1 -: word_length]};
assign pixels_35_19 = {data_out[1280*word_length-1 -: word_length]};
assign pixels_35_20 = {data_out[1281*word_length-1 -: word_length]};
assign pixels_35_21 = {data_out[1282*word_length-1 -: word_length]};
assign pixels_35_22 = {data_out[1283*word_length-1 -: word_length]};
assign pixels_35_23 = {data_out[1284*word_length-1 -: word_length]};
assign pixels_35_24 = {data_out[1285*word_length-1 -: word_length]};
assign pixels_35_25 = {data_out[1286*word_length-1 -: word_length]};
assign pixels_35_26 = {data_out[1287*word_length-1 -: word_length]};
assign pixels_35_27 = {data_out[1288*word_length-1 -: word_length]};
assign pixels_35_28 = {data_out[1289*word_length-1 -: word_length]};
assign pixels_35_29 = {data_out[1290*word_length-1 -: word_length]};
assign pixels_35_30 = {data_out[1291*word_length-1 -: word_length]};
assign pixels_35_31 = {data_out[1292*word_length-1 -: word_length]};
assign pixels_35_32 = {data_out[1293*word_length-1 -: word_length]};
assign pixels_35_33 = {data_out[1294*word_length-1 -: word_length]};
assign pixels_35_34 = {data_out[1295*word_length-1 -: word_length]};
assign pixels_35_35 = {data_out[1296*word_length-1 -: word_length]};

wire [col_length-1:0] pixels_col_0_0, pixels_row_0_0, pixels_col_0_1, pixels_row_0_1, pixels_col_0_2, pixels_row_0_2, pixels_col_0_3, pixels_row_0_3, pixels_col_0_4, pixels_row_0_4, pixels_col_0_5, pixels_row_0_5, pixels_col_0_6, pixels_row_0_6, pixels_col_0_7, pixels_row_0_7, pixels_col_0_8, pixels_row_0_8, pixels_col_0_9, pixels_row_0_9, pixels_col_0_10, pixels_row_0_10, pixels_col_0_11, pixels_row_0_11, pixels_col_0_12, pixels_row_0_12, pixels_col_0_13, pixels_row_0_13, pixels_col_0_14, pixels_row_0_14, pixels_col_0_15, pixels_row_0_15, pixels_col_0_16, pixels_row_0_16, pixels_col_0_17, pixels_row_0_17, pixels_col_0_18, pixels_row_0_18, pixels_col_0_19, pixels_row_0_19, pixels_col_0_20, pixels_row_0_20, pixels_col_0_21, pixels_row_0_21, pixels_col_0_22, pixels_row_0_22, pixels_col_0_23, pixels_row_0_23, pixels_col_0_24, pixels_row_0_24, pixels_col_0_25, pixels_row_0_25, pixels_col_0_26, pixels_row_0_26, pixels_col_0_27, pixels_row_0_27, pixels_col_0_28, pixels_row_0_28, pixels_col_0_29, pixels_row_0_29, pixels_col_0_30, pixels_row_0_30, pixels_col_0_31, pixels_row_0_31, pixels_col_0_32, pixels_row_0_32, pixels_col_0_33, pixels_row_0_33, pixels_col_0_34, pixels_row_0_34, pixels_col_0_35, pixels_row_0_35, pixels_col_1_0, pixels_row_1_0, pixels_col_1_1, pixels_row_1_1, pixels_col_1_2, pixels_row_1_2, pixels_col_1_3, pixels_row_1_3, pixels_col_1_4, pixels_row_1_4, pixels_col_1_5, pixels_row_1_5, pixels_col_1_6, pixels_row_1_6, pixels_col_1_7, pixels_row_1_7, pixels_col_1_8, pixels_row_1_8, pixels_col_1_9, pixels_row_1_9, pixels_col_1_10, pixels_row_1_10, pixels_col_1_11, pixels_row_1_11, pixels_col_1_12, pixels_row_1_12, pixels_col_1_13, pixels_row_1_13, pixels_col_1_14, pixels_row_1_14, pixels_col_1_15, pixels_row_1_15, pixels_col_1_16, pixels_row_1_16, pixels_col_1_17, pixels_row_1_17, pixels_col_1_18, pixels_row_1_18, pixels_col_1_19, pixels_row_1_19, pixels_col_1_20, pixels_row_1_20, pixels_col_1_21, pixels_row_1_21, pixels_col_1_22, pixels_row_1_22, pixels_col_1_23, pixels_row_1_23, pixels_col_1_24, pixels_row_1_24, pixels_col_1_25, pixels_row_1_25, pixels_col_1_26, pixels_row_1_26, pixels_col_1_27, pixels_row_1_27, pixels_col_1_28, pixels_row_1_28, pixels_col_1_29, pixels_row_1_29, pixels_col_1_30, pixels_row_1_30, pixels_col_1_31, pixels_row_1_31, pixels_col_1_32, pixels_row_1_32, pixels_col_1_33, pixels_row_1_33, pixels_col_1_34, pixels_row_1_34, pixels_col_1_35, pixels_row_1_35, pixels_col_2_0, pixels_row_2_0, pixels_col_2_1, pixels_row_2_1, pixels_col_2_2, pixels_row_2_2, pixels_col_2_3, pixels_row_2_3, pixels_col_2_4, pixels_row_2_4, pixels_col_2_5, pixels_row_2_5, pixels_col_2_6, pixels_row_2_6, pixels_col_2_7, pixels_row_2_7, pixels_col_2_8, pixels_row_2_8, pixels_col_2_9, pixels_row_2_9, pixels_col_2_10, pixels_row_2_10, pixels_col_2_11, pixels_row_2_11, pixels_col_2_12, pixels_row_2_12, pixels_col_2_13, pixels_row_2_13, pixels_col_2_14, pixels_row_2_14, pixels_col_2_15, pixels_row_2_15, pixels_col_2_16, pixels_row_2_16, pixels_col_2_17, pixels_row_2_17, pixels_col_2_18, pixels_row_2_18, pixels_col_2_19, pixels_row_2_19, pixels_col_2_20, pixels_row_2_20, pixels_col_2_21, pixels_row_2_21, pixels_col_2_22, pixels_row_2_22, pixels_col_2_23, pixels_row_2_23, pixels_col_2_24, pixels_row_2_24, pixels_col_2_25, pixels_row_2_25, pixels_col_2_26, pixels_row_2_26, pixels_col_2_27, pixels_row_2_27, pixels_col_2_28, pixels_row_2_28, pixels_col_2_29, pixels_row_2_29, pixels_col_2_30, pixels_row_2_30, pixels_col_2_31, pixels_row_2_31, pixels_col_2_32, pixels_row_2_32, pixels_col_2_33, pixels_row_2_33, pixels_col_2_34, pixels_row_2_34, pixels_col_2_35, pixels_row_2_35, pixels_col_3_0, pixels_row_3_0, pixels_col_3_1, pixels_row_3_1, pixels_col_3_2, pixels_row_3_2, pixels_col_3_3, pixels_row_3_3, pixels_col_3_4, pixels_row_3_4, pixels_col_3_5, pixels_row_3_5, pixels_col_3_6, pixels_row_3_6, pixels_col_3_7, pixels_row_3_7, pixels_col_3_8, pixels_row_3_8, pixels_col_3_9, pixels_row_3_9, pixels_col_3_10, pixels_row_3_10, pixels_col_3_11, pixels_row_3_11, pixels_col_3_12, pixels_row_3_12, pixels_col_3_13, pixels_row_3_13, pixels_col_3_14, pixels_row_3_14, pixels_col_3_15, pixels_row_3_15, pixels_col_3_16, pixels_row_3_16, pixels_col_3_17, pixels_row_3_17, pixels_col_3_18, pixels_row_3_18, pixels_col_3_19, pixels_row_3_19, pixels_col_3_20, pixels_row_3_20, pixels_col_3_21, pixels_row_3_21, pixels_col_3_22, pixels_row_3_22, pixels_col_3_23, pixels_row_3_23, pixels_col_3_24, pixels_row_3_24, pixels_col_3_25, pixels_row_3_25, pixels_col_3_26, pixels_row_3_26, pixels_col_3_27, pixels_row_3_27, pixels_col_3_28, pixels_row_3_28, pixels_col_3_29, pixels_row_3_29, pixels_col_3_30, pixels_row_3_30, pixels_col_3_31, pixels_row_3_31, pixels_col_3_32, pixels_row_3_32, pixels_col_3_33, pixels_row_3_33, pixels_col_3_34, pixels_row_3_34, pixels_col_3_35, pixels_row_3_35, pixels_col_4_0, pixels_row_4_0, pixels_col_4_1, pixels_row_4_1, pixels_col_4_2, pixels_row_4_2, pixels_col_4_3, pixels_row_4_3, pixels_col_4_4, pixels_row_4_4, pixels_col_4_5, pixels_row_4_5, pixels_col_4_6, pixels_row_4_6, pixels_col_4_7, pixels_row_4_7, pixels_col_4_8, pixels_row_4_8, pixels_col_4_9, pixels_row_4_9, pixels_col_4_10, pixels_row_4_10, pixels_col_4_11, pixels_row_4_11, pixels_col_4_12, pixels_row_4_12, pixels_col_4_13, pixels_row_4_13, pixels_col_4_14, pixels_row_4_14, pixels_col_4_15, pixels_row_4_15, pixels_col_4_16, pixels_row_4_16, pixels_col_4_17, pixels_row_4_17, pixels_col_4_18, pixels_row_4_18, pixels_col_4_19, pixels_row_4_19, pixels_col_4_20, pixels_row_4_20, pixels_col_4_21, pixels_row_4_21, pixels_col_4_22, pixels_row_4_22, pixels_col_4_23, pixels_row_4_23, pixels_col_4_24, pixels_row_4_24, pixels_col_4_25, pixels_row_4_25, pixels_col_4_26, pixels_row_4_26, pixels_col_4_27, pixels_row_4_27, pixels_col_4_28, pixels_row_4_28, pixels_col_4_29, pixels_row_4_29, pixels_col_4_30, pixels_row_4_30, pixels_col_4_31, pixels_row_4_31, pixels_col_4_32, pixels_row_4_32, pixels_col_4_33, pixels_row_4_33, pixels_col_4_34, pixels_row_4_34, pixels_col_4_35, pixels_row_4_35, pixels_col_5_0, pixels_row_5_0, pixels_col_5_1, pixels_row_5_1, pixels_col_5_2, pixels_row_5_2, pixels_col_5_3, pixels_row_5_3, pixels_col_5_4, pixels_row_5_4, pixels_col_5_5, pixels_row_5_5, pixels_col_5_6, pixels_row_5_6, pixels_col_5_7, pixels_row_5_7, pixels_col_5_8, pixels_row_5_8, pixels_col_5_9, pixels_row_5_9, pixels_col_5_10, pixels_row_5_10, pixels_col_5_11, pixels_row_5_11, pixels_col_5_12, pixels_row_5_12, pixels_col_5_13, pixels_row_5_13, pixels_col_5_14, pixels_row_5_14, pixels_col_5_15, pixels_row_5_15, pixels_col_5_16, pixels_row_5_16, pixels_col_5_17, pixels_row_5_17, pixels_col_5_18, pixels_row_5_18, pixels_col_5_19, pixels_row_5_19, pixels_col_5_20, pixels_row_5_20, pixels_col_5_21, pixels_row_5_21, pixels_col_5_22, pixels_row_5_22, pixels_col_5_23, pixels_row_5_23, pixels_col_5_24, pixels_row_5_24, pixels_col_5_25, pixels_row_5_25, pixels_col_5_26, pixels_row_5_26, pixels_col_5_27, pixels_row_5_27, pixels_col_5_28, pixels_row_5_28, pixels_col_5_29, pixels_row_5_29, pixels_col_5_30, pixels_row_5_30, pixels_col_5_31, pixels_row_5_31, pixels_col_5_32, pixels_row_5_32, pixels_col_5_33, pixels_row_5_33, pixels_col_5_34, pixels_row_5_34, pixels_col_5_35, pixels_row_5_35, pixels_col_6_0, pixels_row_6_0, pixels_col_6_1, pixels_row_6_1, pixels_col_6_2, pixels_row_6_2, pixels_col_6_3, pixels_row_6_3, pixels_col_6_4, pixels_row_6_4, pixels_col_6_5, pixels_row_6_5, pixels_col_6_6, pixels_row_6_6, pixels_col_6_7, pixels_row_6_7, pixels_col_6_8, pixels_row_6_8, pixels_col_6_9, pixels_row_6_9, pixels_col_6_10, pixels_row_6_10, pixels_col_6_11, pixels_row_6_11, pixels_col_6_12, pixels_row_6_12, pixels_col_6_13, pixels_row_6_13, pixels_col_6_14, pixels_row_6_14, pixels_col_6_15, pixels_row_6_15, pixels_col_6_16, pixels_row_6_16, pixels_col_6_17, pixels_row_6_17, pixels_col_6_18, pixels_row_6_18, pixels_col_6_19, pixels_row_6_19, pixels_col_6_20, pixels_row_6_20, pixels_col_6_21, pixels_row_6_21, pixels_col_6_22, pixels_row_6_22, pixels_col_6_23, pixels_row_6_23, pixels_col_6_24, pixels_row_6_24, pixels_col_6_25, pixels_row_6_25, pixels_col_6_26, pixels_row_6_26, pixels_col_6_27, pixels_row_6_27, pixels_col_6_28, pixels_row_6_28, pixels_col_6_29, pixels_row_6_29, pixels_col_6_30, pixels_row_6_30, pixels_col_6_31, pixels_row_6_31, pixels_col_6_32, pixels_row_6_32, pixels_col_6_33, pixels_row_6_33, pixels_col_6_34, pixels_row_6_34, pixels_col_6_35, pixels_row_6_35, pixels_col_7_0, pixels_row_7_0, pixels_col_7_1, pixels_row_7_1, pixels_col_7_2, pixels_row_7_2, pixels_col_7_3, pixels_row_7_3, pixels_col_7_4, pixels_row_7_4, pixels_col_7_5, pixels_row_7_5, pixels_col_7_6, pixels_row_7_6, pixels_col_7_7, pixels_row_7_7, pixels_col_7_8, pixels_row_7_8, pixels_col_7_9, pixels_row_7_9, pixels_col_7_10, pixels_row_7_10, pixels_col_7_11, pixels_row_7_11, pixels_col_7_12, pixels_row_7_12, pixels_col_7_13, pixels_row_7_13, pixels_col_7_14, pixels_row_7_14, pixels_col_7_15, pixels_row_7_15, pixels_col_7_16, pixels_row_7_16, pixels_col_7_17, pixels_row_7_17, pixels_col_7_18, pixels_row_7_18, pixels_col_7_19, pixels_row_7_19, pixels_col_7_20, pixels_row_7_20, pixels_col_7_21, pixels_row_7_21, pixels_col_7_22, pixels_row_7_22, pixels_col_7_23, pixels_row_7_23, pixels_col_7_24, pixels_row_7_24, pixels_col_7_25, pixels_row_7_25, pixels_col_7_26, pixels_row_7_26, pixels_col_7_27, pixels_row_7_27, pixels_col_7_28, pixels_row_7_28, pixels_col_7_29, pixels_row_7_29, pixels_col_7_30, pixels_row_7_30, pixels_col_7_31, pixels_row_7_31, pixels_col_7_32, pixels_row_7_32, pixels_col_7_33, pixels_row_7_33, pixels_col_7_34, pixels_row_7_34, pixels_col_7_35, pixels_row_7_35, pixels_col_8_0, pixels_row_8_0, pixels_col_8_1, pixels_row_8_1, pixels_col_8_2, pixels_row_8_2, pixels_col_8_3, pixels_row_8_3, pixels_col_8_4, pixels_row_8_4, pixels_col_8_5, pixels_row_8_5, pixels_col_8_6, pixels_row_8_6, pixels_col_8_7, pixels_row_8_7, pixels_col_8_8, pixels_row_8_8, pixels_col_8_9, pixels_row_8_9, 
pixels_col_8_10, pixels_row_8_10, pixels_col_8_11, pixels_row_8_11, pixels_col_8_12, pixels_row_8_12, pixels_col_8_13, pixels_row_8_13, pixels_col_8_14, pixels_row_8_14, pixels_col_8_15, pixels_row_8_15, pixels_col_8_16, pixels_row_8_16, pixels_col_8_17, pixels_row_8_17, pixels_col_8_18, pixels_row_8_18, pixels_col_8_19, pixels_row_8_19, pixels_col_8_20, pixels_row_8_20, pixels_col_8_21, pixels_row_8_21, pixels_col_8_22, pixels_row_8_22, pixels_col_8_23, pixels_row_8_23, pixels_col_8_24, pixels_row_8_24, pixels_col_8_25, pixels_row_8_25, pixels_col_8_26, pixels_row_8_26, pixels_col_8_27, pixels_row_8_27, pixels_col_8_28, pixels_row_8_28, pixels_col_8_29, pixels_row_8_29, pixels_col_8_30, pixels_row_8_30, pixels_col_8_31, pixels_row_8_31, pixels_col_8_32, pixels_row_8_32, pixels_col_8_33, pixels_row_8_33, pixels_col_8_34, pixels_row_8_34, pixels_col_8_35, pixels_row_8_35, pixels_col_9_0, pixels_row_9_0, pixels_col_9_1, pixels_row_9_1, pixels_col_9_2, pixels_row_9_2, pixels_col_9_3, pixels_row_9_3, pixels_col_9_4, pixels_row_9_4, pixels_col_9_5, pixels_row_9_5, pixels_col_9_6, pixels_row_9_6, pixels_col_9_7, pixels_row_9_7, pixels_col_9_8, pixels_row_9_8, pixels_col_9_9, pixels_row_9_9, pixels_col_9_10, pixels_row_9_10, pixels_col_9_11, pixels_row_9_11, pixels_col_9_12, pixels_row_9_12, pixels_col_9_13, pixels_row_9_13, pixels_col_9_14, pixels_row_9_14, pixels_col_9_15, pixels_row_9_15, pixels_col_9_16, pixels_row_9_16, pixels_col_9_17, pixels_row_9_17, pixels_col_9_18, pixels_row_9_18, pixels_col_9_19, pixels_row_9_19, pixels_col_9_20, pixels_row_9_20, pixels_col_9_21, pixels_row_9_21, pixels_col_9_22, pixels_row_9_22, pixels_col_9_23, pixels_row_9_23, pixels_col_9_24, pixels_row_9_24, pixels_col_9_25, pixels_row_9_25, pixels_col_9_26, pixels_row_9_26, pixels_col_9_27, pixels_row_9_27, pixels_col_9_28, pixels_row_9_28, pixels_col_9_29, pixels_row_9_29, pixels_col_9_30, pixels_row_9_30, pixels_col_9_31, pixels_row_9_31, pixels_col_9_32, pixels_row_9_32, pixels_col_9_33, pixels_row_9_33, pixels_col_9_34, pixels_row_9_34, pixels_col_9_35, pixels_row_9_35, pixels_col_10_0, pixels_row_10_0, pixels_col_10_1, pixels_row_10_1, pixels_col_10_2, pixels_row_10_2, pixels_col_10_3, pixels_row_10_3, pixels_col_10_4, pixels_row_10_4, pixels_col_10_5, pixels_row_10_5, pixels_col_10_6, pixels_row_10_6, pixels_col_10_7, pixels_row_10_7, pixels_col_10_8, pixels_row_10_8, pixels_col_10_9, pixels_row_10_9, pixels_col_10_10, pixels_row_10_10, pixels_col_10_11, pixels_row_10_11, pixels_col_10_12, pixels_row_10_12, pixels_col_10_13, pixels_row_10_13, pixels_col_10_14, pixels_row_10_14, pixels_col_10_15, pixels_row_10_15, pixels_col_10_16, pixels_row_10_16, pixels_col_10_17, pixels_row_10_17, pixels_col_10_18, pixels_row_10_18, pixels_col_10_19, pixels_row_10_19, pixels_col_10_20, pixels_row_10_20, pixels_col_10_21, pixels_row_10_21, pixels_col_10_22, pixels_row_10_22, pixels_col_10_23, pixels_row_10_23, pixels_col_10_24, pixels_row_10_24, pixels_col_10_25, pixels_row_10_25, pixels_col_10_26, pixels_row_10_26, pixels_col_10_27, pixels_row_10_27, pixels_col_10_28, pixels_row_10_28, pixels_col_10_29, pixels_row_10_29, pixels_col_10_30, pixels_row_10_30, pixels_col_10_31, pixels_row_10_31, pixels_col_10_32, pixels_row_10_32, pixels_col_10_33, pixels_row_10_33, pixels_col_10_34, pixels_row_10_34, pixels_col_10_35, pixels_row_10_35, pixels_col_11_0, pixels_row_11_0, pixels_col_11_1, pixels_row_11_1, pixels_col_11_2, pixels_row_11_2, pixels_col_11_3, pixels_row_11_3, pixels_col_11_4, pixels_row_11_4, pixels_col_11_5, pixels_row_11_5, pixels_col_11_6, pixels_row_11_6, pixels_col_11_7, pixels_row_11_7, pixels_col_11_8, pixels_row_11_8, pixels_col_11_9, pixels_row_11_9, pixels_col_11_10, pixels_row_11_10, pixels_col_11_11, pixels_row_11_11, pixels_col_11_12, pixels_row_11_12, pixels_col_11_13, pixels_row_11_13, pixels_col_11_14, pixels_row_11_14, pixels_col_11_15, pixels_row_11_15, pixels_col_11_16, pixels_row_11_16, pixels_col_11_17, pixels_row_11_17, pixels_col_11_18, pixels_row_11_18, pixels_col_11_19, pixels_row_11_19, pixels_col_11_20, pixels_row_11_20, pixels_col_11_21, pixels_row_11_21, pixels_col_11_22, pixels_row_11_22, pixels_col_11_23, pixels_row_11_23, pixels_col_11_24, pixels_row_11_24, pixels_col_11_25, pixels_row_11_25, pixels_col_11_26, pixels_row_11_26, pixels_col_11_27, pixels_row_11_27, pixels_col_11_28, pixels_row_11_28, pixels_col_11_29, pixels_row_11_29, pixels_col_11_30, pixels_row_11_30, pixels_col_11_31, pixels_row_11_31, pixels_col_11_32, pixels_row_11_32, pixels_col_11_33, pixels_row_11_33, pixels_col_11_34, pixels_row_11_34, pixels_col_11_35, pixels_row_11_35, pixels_col_12_0, pixels_row_12_0, pixels_col_12_1, pixels_row_12_1, pixels_col_12_2, pixels_row_12_2, pixels_col_12_3, pixels_row_12_3, pixels_col_12_4, pixels_row_12_4, pixels_col_12_5, pixels_row_12_5, pixels_col_12_6, pixels_row_12_6, pixels_col_12_7, pixels_row_12_7, pixels_col_12_8, pixels_row_12_8, pixels_col_12_9, pixels_row_12_9, pixels_col_12_10, pixels_row_12_10, pixels_col_12_11, pixels_row_12_11, pixels_col_12_12, pixels_row_12_12, pixels_col_12_13, pixels_row_12_13, pixels_col_12_14, pixels_row_12_14, pixels_col_12_15, pixels_row_12_15, pixels_col_12_16, pixels_row_12_16, pixels_col_12_17, pixels_row_12_17, pixels_col_12_18, pixels_row_12_18, pixels_col_12_19, pixels_row_12_19, pixels_col_12_20, pixels_row_12_20, pixels_col_12_21, pixels_row_12_21, pixels_col_12_22, pixels_row_12_22, pixels_col_12_23, pixels_row_12_23, pixels_col_12_24, pixels_row_12_24, pixels_col_12_25, pixels_row_12_25, pixels_col_12_26, pixels_row_12_26, pixels_col_12_27, pixels_row_12_27, pixels_col_12_28, pixels_row_12_28, pixels_col_12_29, pixels_row_12_29, pixels_col_12_30, pixels_row_12_30, pixels_col_12_31, pixels_row_12_31, pixels_col_12_32, pixels_row_12_32, pixels_col_12_33, pixels_row_12_33, pixels_col_12_34, pixels_row_12_34, pixels_col_12_35, pixels_row_12_35, pixels_col_13_0, pixels_row_13_0, pixels_col_13_1, pixels_row_13_1, pixels_col_13_2, pixels_row_13_2, pixels_col_13_3, pixels_row_13_3, pixels_col_13_4, pixels_row_13_4, pixels_col_13_5, pixels_row_13_5, pixels_col_13_6, pixels_row_13_6, pixels_col_13_7, pixels_row_13_7, pixels_col_13_8, pixels_row_13_8, pixels_col_13_9, pixels_row_13_9, pixels_col_13_10, pixels_row_13_10, pixels_col_13_11, pixels_row_13_11, pixels_col_13_12, pixels_row_13_12, pixels_col_13_13, pixels_row_13_13, pixels_col_13_14, pixels_row_13_14, pixels_col_13_15, pixels_row_13_15, pixels_col_13_16, pixels_row_13_16, pixels_col_13_17, pixels_row_13_17, pixels_col_13_18, pixels_row_13_18, pixels_col_13_19, pixels_row_13_19, pixels_col_13_20, pixels_row_13_20, pixels_col_13_21, pixels_row_13_21, pixels_col_13_22, pixels_row_13_22, pixels_col_13_23, pixels_row_13_23, pixels_col_13_24, pixels_row_13_24, pixels_col_13_25, pixels_row_13_25, pixels_col_13_26, pixels_row_13_26, pixels_col_13_27, pixels_row_13_27, pixels_col_13_28, pixels_row_13_28, pixels_col_13_29, pixels_row_13_29, pixels_col_13_30, pixels_row_13_30, pixels_col_13_31, pixels_row_13_31, pixels_col_13_32, pixels_row_13_32, pixels_col_13_33, pixels_row_13_33, pixels_col_13_34, pixels_row_13_34, pixels_col_13_35, pixels_row_13_35, pixels_col_14_0, pixels_row_14_0, pixels_col_14_1, pixels_row_14_1, pixels_col_14_2, pixels_row_14_2, pixels_col_14_3, pixels_row_14_3, pixels_col_14_4, pixels_row_14_4, pixels_col_14_5, pixels_row_14_5, pixels_col_14_6, pixels_row_14_6, pixels_col_14_7, pixels_row_14_7, pixels_col_14_8, pixels_row_14_8, pixels_col_14_9, pixels_row_14_9, pixels_col_14_10, pixels_row_14_10, pixels_col_14_11, pixels_row_14_11, pixels_col_14_12, pixels_row_14_12, pixels_col_14_13, pixels_row_14_13, pixels_col_14_14, pixels_row_14_14, pixels_col_14_15, pixels_row_14_15, pixels_col_14_16, pixels_row_14_16, pixels_col_14_17, pixels_row_14_17, pixels_col_14_18, pixels_row_14_18, pixels_col_14_19, pixels_row_14_19, pixels_col_14_20, pixels_row_14_20, pixels_col_14_21, pixels_row_14_21, pixels_col_14_22, pixels_row_14_22, pixels_col_14_23, pixels_row_14_23, pixels_col_14_24, pixels_row_14_24, pixels_col_14_25, pixels_row_14_25, pixels_col_14_26, pixels_row_14_26, pixels_col_14_27, pixels_row_14_27, pixels_col_14_28, pixels_row_14_28, pixels_col_14_29, pixels_row_14_29, pixels_col_14_30, pixels_row_14_30, pixels_col_14_31, pixels_row_14_31, pixels_col_14_32, pixels_row_14_32, pixels_col_14_33, pixels_row_14_33, pixels_col_14_34, pixels_row_14_34, pixels_col_14_35, pixels_row_14_35, pixels_col_15_0, pixels_row_15_0, pixels_col_15_1, pixels_row_15_1, pixels_col_15_2, pixels_row_15_2, pixels_col_15_3, pixels_row_15_3, pixels_col_15_4, pixels_row_15_4, pixels_col_15_5, pixels_row_15_5, pixels_col_15_6, pixels_row_15_6, pixels_col_15_7, pixels_row_15_7, pixels_col_15_8, pixels_row_15_8, pixels_col_15_9, pixels_row_15_9, pixels_col_15_10, pixels_row_15_10, pixels_col_15_11, pixels_row_15_11, pixels_col_15_12, pixels_row_15_12, pixels_col_15_13, pixels_row_15_13, pixels_col_15_14, pixels_row_15_14, pixels_col_15_15, pixels_row_15_15, pixels_col_15_16, pixels_row_15_16, pixels_col_15_17, pixels_row_15_17, pixels_col_15_18, pixels_row_15_18, pixels_col_15_19, pixels_row_15_19, pixels_col_15_20, pixels_row_15_20, pixels_col_15_21, pixels_row_15_21, pixels_col_15_22, pixels_row_15_22, pixels_col_15_23, pixels_row_15_23, pixels_col_15_24, pixels_row_15_24, pixels_col_15_25, pixels_row_15_25, pixels_col_15_26, pixels_row_15_26, pixels_col_15_27, pixels_row_15_27, pixels_col_15_28, pixels_row_15_28, pixels_col_15_29, pixels_row_15_29, pixels_col_15_30, pixels_row_15_30, pixels_col_15_31, pixels_row_15_31, pixels_col_15_32, pixels_row_15_32, pixels_col_15_33, pixels_row_15_33, pixels_col_15_34, pixels_row_15_34, pixels_col_15_35, pixels_row_15_35, pixels_col_16_0, pixels_row_16_0, pixels_col_16_1, pixels_row_16_1, pixels_col_16_2, pixels_row_16_2, pixels_col_16_3, pixels_row_16_3, pixels_col_16_4, pixels_row_16_4, pixels_col_16_5, pixels_row_16_5, pixels_col_16_6, pixels_row_16_6, 
pixels_col_16_7, pixels_row_16_7, pixels_col_16_8, pixels_row_16_8, pixels_col_16_9, pixels_row_16_9, pixels_col_16_10, pixels_row_16_10, pixels_col_16_11, pixels_row_16_11, pixels_col_16_12, pixels_row_16_12, pixels_col_16_13, pixels_row_16_13, pixels_col_16_14, pixels_row_16_14, pixels_col_16_15, pixels_row_16_15, pixels_col_16_16, pixels_row_16_16, pixels_col_16_17, pixels_row_16_17, pixels_col_16_18, pixels_row_16_18, pixels_col_16_19, pixels_row_16_19, pixels_col_16_20, pixels_row_16_20, pixels_col_16_21, pixels_row_16_21, pixels_col_16_22, pixels_row_16_22, pixels_col_16_23, pixels_row_16_23, pixels_col_16_24, pixels_row_16_24, pixels_col_16_25, pixels_row_16_25, pixels_col_16_26, pixels_row_16_26, pixels_col_16_27, pixels_row_16_27, pixels_col_16_28, pixels_row_16_28, pixels_col_16_29, pixels_row_16_29, pixels_col_16_30, pixels_row_16_30, pixels_col_16_31, pixels_row_16_31, pixels_col_16_32, pixels_row_16_32, pixels_col_16_33, pixels_row_16_33, pixels_col_16_34, pixels_row_16_34, pixels_col_16_35, pixels_row_16_35, pixels_col_17_0, pixels_row_17_0, pixels_col_17_1, pixels_row_17_1, pixels_col_17_2, pixels_row_17_2, pixels_col_17_3, pixels_row_17_3, pixels_col_17_4, pixels_row_17_4, pixels_col_17_5, pixels_row_17_5, pixels_col_17_6, pixels_row_17_6, pixels_col_17_7, pixels_row_17_7, pixels_col_17_8, pixels_row_17_8, pixels_col_17_9, pixels_row_17_9, pixels_col_17_10, pixels_row_17_10, pixels_col_17_11, pixels_row_17_11, pixels_col_17_12, pixels_row_17_12, pixels_col_17_13, pixels_row_17_13, pixels_col_17_14, pixels_row_17_14, pixels_col_17_15, pixels_row_17_15, pixels_col_17_16, pixels_row_17_16, pixels_col_17_17, pixels_row_17_17, pixels_col_17_18, pixels_row_17_18, pixels_col_17_19, pixels_row_17_19, pixels_col_17_20, pixels_row_17_20, pixels_col_17_21, pixels_row_17_21, pixels_col_17_22, pixels_row_17_22, pixels_col_17_23, pixels_row_17_23, pixels_col_17_24, pixels_row_17_24, pixels_col_17_25, pixels_row_17_25, pixels_col_17_26, pixels_row_17_26, pixels_col_17_27, pixels_row_17_27, pixels_col_17_28, pixels_row_17_28, pixels_col_17_29, pixels_row_17_29, pixels_col_17_30, pixels_row_17_30, pixels_col_17_31, pixels_row_17_31, pixels_col_17_32, pixels_row_17_32, pixels_col_17_33, pixels_row_17_33, pixels_col_17_34, pixels_row_17_34, pixels_col_17_35, pixels_row_17_35, pixels_col_18_0, pixels_row_18_0, pixels_col_18_1, pixels_row_18_1, pixels_col_18_2, pixels_row_18_2, pixels_col_18_3, pixels_row_18_3, pixels_col_18_4, pixels_row_18_4, pixels_col_18_5, pixels_row_18_5, pixels_col_18_6, pixels_row_18_6, pixels_col_18_7, pixels_row_18_7, pixels_col_18_8, pixels_row_18_8, pixels_col_18_9, pixels_row_18_9, pixels_col_18_10, pixels_row_18_10, pixels_col_18_11, pixels_row_18_11, pixels_col_18_12, pixels_row_18_12, pixels_col_18_13, pixels_row_18_13, pixels_col_18_14, pixels_row_18_14, pixels_col_18_15, pixels_row_18_15, pixels_col_18_16, pixels_row_18_16, pixels_col_18_17, pixels_row_18_17, pixels_col_18_18, pixels_row_18_18, pixels_col_18_19, pixels_row_18_19, pixels_col_18_20, pixels_row_18_20, pixels_col_18_21, pixels_row_18_21, pixels_col_18_22, pixels_row_18_22, pixels_col_18_23, pixels_row_18_23, pixels_col_18_24, pixels_row_18_24, pixels_col_18_25, pixels_row_18_25, pixels_col_18_26, pixels_row_18_26, pixels_col_18_27, pixels_row_18_27, pixels_col_18_28, pixels_row_18_28, pixels_col_18_29, pixels_row_18_29, pixels_col_18_30, pixels_row_18_30, pixels_col_18_31, pixels_row_18_31, pixels_col_18_32, pixels_row_18_32, pixels_col_18_33, pixels_row_18_33, pixels_col_18_34, pixels_row_18_34, pixels_col_18_35, pixels_row_18_35, pixels_col_19_0, pixels_row_19_0, pixels_col_19_1, pixels_row_19_1, pixels_col_19_2, pixels_row_19_2, pixels_col_19_3, pixels_row_19_3, pixels_col_19_4, pixels_row_19_4, pixels_col_19_5, pixels_row_19_5, pixels_col_19_6, pixels_row_19_6, pixels_col_19_7, pixels_row_19_7, pixels_col_19_8, pixels_row_19_8, pixels_col_19_9, pixels_row_19_9, pixels_col_19_10, pixels_row_19_10, pixels_col_19_11, pixels_row_19_11, pixels_col_19_12, pixels_row_19_12, pixels_col_19_13, pixels_row_19_13, pixels_col_19_14, pixels_row_19_14, pixels_col_19_15, pixels_row_19_15, pixels_col_19_16, pixels_row_19_16, pixels_col_19_17, pixels_row_19_17, pixels_col_19_18, pixels_row_19_18, pixels_col_19_19, pixels_row_19_19, pixels_col_19_20, pixels_row_19_20, pixels_col_19_21, pixels_row_19_21, pixels_col_19_22, pixels_row_19_22, pixels_col_19_23, pixels_row_19_23, pixels_col_19_24, pixels_row_19_24, pixels_col_19_25, pixels_row_19_25, pixels_col_19_26, pixels_row_19_26, pixels_col_19_27, pixels_row_19_27, pixels_col_19_28, pixels_row_19_28, pixels_col_19_29, pixels_row_19_29, pixels_col_19_30, pixels_row_19_30, pixels_col_19_31, pixels_row_19_31, pixels_col_19_32, pixels_row_19_32, pixels_col_19_33, pixels_row_19_33, pixels_col_19_34, pixels_row_19_34, pixels_col_19_35, pixels_row_19_35, pixels_col_20_0, pixels_row_20_0, pixels_col_20_1, pixels_row_20_1, pixels_col_20_2, pixels_row_20_2, pixels_col_20_3, pixels_row_20_3, pixels_col_20_4, pixels_row_20_4, pixels_col_20_5, pixels_row_20_5, pixels_col_20_6, pixels_row_20_6, pixels_col_20_7, pixels_row_20_7, pixels_col_20_8, pixels_row_20_8, pixels_col_20_9, pixels_row_20_9, pixels_col_20_10, pixels_row_20_10, pixels_col_20_11, pixels_row_20_11, pixels_col_20_12, pixels_row_20_12, pixels_col_20_13, pixels_row_20_13, pixels_col_20_14, pixels_row_20_14, pixels_col_20_15, pixels_row_20_15, pixels_col_20_16, pixels_row_20_16, pixels_col_20_17, pixels_row_20_17, pixels_col_20_18, pixels_row_20_18, pixels_col_20_19, pixels_row_20_19, pixels_col_20_20, pixels_row_20_20, pixels_col_20_21, pixels_row_20_21, pixels_col_20_22, pixels_row_20_22, pixels_col_20_23, pixels_row_20_23, pixels_col_20_24, pixels_row_20_24, pixels_col_20_25, pixels_row_20_25, pixels_col_20_26, pixels_row_20_26, pixels_col_20_27, pixels_row_20_27, pixels_col_20_28, pixels_row_20_28, pixels_col_20_29, pixels_row_20_29, pixels_col_20_30, pixels_row_20_30, pixels_col_20_31, pixels_row_20_31, pixels_col_20_32, pixels_row_20_32, pixels_col_20_33, pixels_row_20_33, pixels_col_20_34, pixels_row_20_34, pixels_col_20_35, pixels_row_20_35, pixels_col_21_0, pixels_row_21_0, pixels_col_21_1, pixels_row_21_1, pixels_col_21_2, pixels_row_21_2, pixels_col_21_3, pixels_row_21_3, pixels_col_21_4, pixels_row_21_4, pixels_col_21_5, pixels_row_21_5, pixels_col_21_6, pixels_row_21_6, pixels_col_21_7, pixels_row_21_7, pixels_col_21_8, pixels_row_21_8, pixels_col_21_9, pixels_row_21_9, pixels_col_21_10, pixels_row_21_10, pixels_col_21_11, pixels_row_21_11, pixels_col_21_12, pixels_row_21_12, pixels_col_21_13, pixels_row_21_13, pixels_col_21_14, pixels_row_21_14, pixels_col_21_15, pixels_row_21_15, pixels_col_21_16, pixels_row_21_16, pixels_col_21_17, pixels_row_21_17, pixels_col_21_18, pixels_row_21_18, pixels_col_21_19, pixels_row_21_19, pixels_col_21_20, pixels_row_21_20, pixels_col_21_21, pixels_row_21_21, pixels_col_21_22, pixels_row_21_22, pixels_col_21_23, pixels_row_21_23, pixels_col_21_24, pixels_row_21_24, pixels_col_21_25, pixels_row_21_25, pixels_col_21_26, pixels_row_21_26, pixels_col_21_27, pixels_row_21_27, pixels_col_21_28, pixels_row_21_28, pixels_col_21_29, pixels_row_21_29, pixels_col_21_30, pixels_row_21_30, pixels_col_21_31, pixels_row_21_31, pixels_col_21_32, pixels_row_21_32, pixels_col_21_33, pixels_row_21_33, pixels_col_21_34, pixels_row_21_34, pixels_col_21_35, pixels_row_21_35, pixels_col_22_0, pixels_row_22_0, pixels_col_22_1, pixels_row_22_1, pixels_col_22_2, pixels_row_22_2, pixels_col_22_3, pixels_row_22_3, pixels_col_22_4, pixels_row_22_4, pixels_col_22_5, pixels_row_22_5, pixels_col_22_6, pixels_row_22_6, pixels_col_22_7, pixels_row_22_7, pixels_col_22_8, pixels_row_22_8, pixels_col_22_9, pixels_row_22_9, pixels_col_22_10, pixels_row_22_10, pixels_col_22_11, pixels_row_22_11, pixels_col_22_12, pixels_row_22_12, pixels_col_22_13, pixels_row_22_13, pixels_col_22_14, pixels_row_22_14, pixels_col_22_15, pixels_row_22_15, pixels_col_22_16, pixels_row_22_16, pixels_col_22_17, pixels_row_22_17, pixels_col_22_18, pixels_row_22_18, pixels_col_22_19, pixels_row_22_19, pixels_col_22_20, pixels_row_22_20, pixels_col_22_21, pixels_row_22_21, pixels_col_22_22, pixels_row_22_22, pixels_col_22_23, pixels_row_22_23, pixels_col_22_24, pixels_row_22_24, pixels_col_22_25, pixels_row_22_25, pixels_col_22_26, pixels_row_22_26, pixels_col_22_27, pixels_row_22_27, pixels_col_22_28, pixels_row_22_28, pixels_col_22_29, pixels_row_22_29, pixels_col_22_30, pixels_row_22_30, pixels_col_22_31, pixels_row_22_31, pixels_col_22_32, pixels_row_22_32, pixels_col_22_33, pixels_row_22_33, pixels_col_22_34, pixels_row_22_34, pixels_col_22_35, pixels_row_22_35, pixels_col_23_0, pixels_row_23_0, pixels_col_23_1, pixels_row_23_1, pixels_col_23_2, pixels_row_23_2, pixels_col_23_3, pixels_row_23_3, pixels_col_23_4, pixels_row_23_4, pixels_col_23_5, pixels_row_23_5, pixels_col_23_6, pixels_row_23_6, pixels_col_23_7, pixels_row_23_7, pixels_col_23_8, pixels_row_23_8, pixels_col_23_9, pixels_row_23_9, pixels_col_23_10, pixels_row_23_10, pixels_col_23_11, pixels_row_23_11, pixels_col_23_12, pixels_row_23_12, pixels_col_23_13, pixels_row_23_13, pixels_col_23_14, pixels_row_23_14, pixels_col_23_15, pixels_row_23_15, pixels_col_23_16, pixels_row_23_16, pixels_col_23_17, pixels_row_23_17, pixels_col_23_18, pixels_row_23_18, pixels_col_23_19, pixels_row_23_19, pixels_col_23_20, pixels_row_23_20, pixels_col_23_21, pixels_row_23_21, pixels_col_23_22, pixels_row_23_22, pixels_col_23_23, pixels_row_23_23, pixels_col_23_24, pixels_row_23_24, pixels_col_23_25, pixels_row_23_25, pixels_col_23_26, pixels_row_23_26, pixels_col_23_27, pixels_row_23_27, pixels_col_23_28, pixels_row_23_28, pixels_col_23_29, pixels_row_23_29, pixels_col_23_30, pixels_row_23_30, pixels_col_23_31, pixels_row_23_31, pixels_col_23_32, pixels_row_23_32, pixels_col_23_33, pixels_row_23_33, pixels_col_23_34, pixels_row_23_34, pixels_col_23_35, pixels_row_23_35, pixels_col_24_0, 
pixels_row_24_0, pixels_col_24_1, pixels_row_24_1, pixels_col_24_2, pixels_row_24_2, pixels_col_24_3, pixels_row_24_3, pixels_col_24_4, pixels_row_24_4, pixels_col_24_5, pixels_row_24_5, pixels_col_24_6, pixels_row_24_6, pixels_col_24_7, pixels_row_24_7, pixels_col_24_8, pixels_row_24_8, pixels_col_24_9, pixels_row_24_9, pixels_col_24_10, pixels_row_24_10, pixels_col_24_11, pixels_row_24_11, pixels_col_24_12, pixels_row_24_12, pixels_col_24_13, pixels_row_24_13, pixels_col_24_14, pixels_row_24_14, pixels_col_24_15, pixels_row_24_15, pixels_col_24_16, pixels_row_24_16, pixels_col_24_17, pixels_row_24_17, pixels_col_24_18, pixels_row_24_18, pixels_col_24_19, pixels_row_24_19, pixels_col_24_20, pixels_row_24_20, pixels_col_24_21, pixels_row_24_21, pixels_col_24_22, pixels_row_24_22, pixels_col_24_23, pixels_row_24_23, pixels_col_24_24, pixels_row_24_24, pixels_col_24_25, pixels_row_24_25, pixels_col_24_26, pixels_row_24_26, pixels_col_24_27, pixels_row_24_27, pixels_col_24_28, pixels_row_24_28, pixels_col_24_29, pixels_row_24_29, pixels_col_24_30, pixels_row_24_30, pixels_col_24_31, pixels_row_24_31, pixels_col_24_32, pixels_row_24_32, pixels_col_24_33, pixels_row_24_33, pixels_col_24_34, pixels_row_24_34, pixels_col_24_35, pixels_row_24_35, pixels_col_25_0, pixels_row_25_0, pixels_col_25_1, pixels_row_25_1, pixels_col_25_2, pixels_row_25_2, pixels_col_25_3, pixels_row_25_3, pixels_col_25_4, pixels_row_25_4, pixels_col_25_5, pixels_row_25_5, pixels_col_25_6, pixels_row_25_6, pixels_col_25_7, pixels_row_25_7, pixels_col_25_8, pixels_row_25_8, pixels_col_25_9, pixels_row_25_9, pixels_col_25_10, pixels_row_25_10, pixels_col_25_11, pixels_row_25_11, pixels_col_25_12, pixels_row_25_12, pixels_col_25_13, pixels_row_25_13, pixels_col_25_14, pixels_row_25_14, pixels_col_25_15, pixels_row_25_15, pixels_col_25_16, pixels_row_25_16, pixels_col_25_17, pixels_row_25_17, pixels_col_25_18, pixels_row_25_18, pixels_col_25_19, pixels_row_25_19, pixels_col_25_20, pixels_row_25_20, pixels_col_25_21, pixels_row_25_21, pixels_col_25_22, pixels_row_25_22, pixels_col_25_23, pixels_row_25_23, pixels_col_25_24, pixels_row_25_24, pixels_col_25_25, pixels_row_25_25, pixels_col_25_26, pixels_row_25_26, pixels_col_25_27, pixels_row_25_27, pixels_col_25_28, pixels_row_25_28, pixels_col_25_29, pixels_row_25_29, pixels_col_25_30, pixels_row_25_30, pixels_col_25_31, pixels_row_25_31, pixels_col_25_32, pixels_row_25_32, pixels_col_25_33, pixels_row_25_33, pixels_col_25_34, pixels_row_25_34, pixels_col_25_35, pixels_row_25_35, pixels_col_26_0, pixels_row_26_0, pixels_col_26_1, pixels_row_26_1, pixels_col_26_2, pixels_row_26_2, pixels_col_26_3, pixels_row_26_3, pixels_col_26_4, pixels_row_26_4, pixels_col_26_5, pixels_row_26_5, pixels_col_26_6, pixels_row_26_6, pixels_col_26_7, pixels_row_26_7, pixels_col_26_8, pixels_row_26_8, pixels_col_26_9, pixels_row_26_9, pixels_col_26_10, pixels_row_26_10, pixels_col_26_11, pixels_row_26_11, pixels_col_26_12, pixels_row_26_12, pixels_col_26_13, pixels_row_26_13, pixels_col_26_14, pixels_row_26_14, pixels_col_26_15, pixels_row_26_15, pixels_col_26_16, pixels_row_26_16, pixels_col_26_17, pixels_row_26_17, pixels_col_26_18, pixels_row_26_18, pixels_col_26_19, pixels_row_26_19, pixels_col_26_20, pixels_row_26_20, pixels_col_26_21, pixels_row_26_21, pixels_col_26_22, pixels_row_26_22, pixels_col_26_23, pixels_row_26_23, pixels_col_26_24, pixels_row_26_24, pixels_col_26_25, pixels_row_26_25, pixels_col_26_26, pixels_row_26_26, pixels_col_26_27, pixels_row_26_27, pixels_col_26_28, pixels_row_26_28, pixels_col_26_29, pixels_row_26_29, pixels_col_26_30, pixels_row_26_30, pixels_col_26_31, pixels_row_26_31, pixels_col_26_32, pixels_row_26_32, pixels_col_26_33, pixels_row_26_33, pixels_col_26_34, pixels_row_26_34, pixels_col_26_35, pixels_row_26_35, pixels_col_27_0, pixels_row_27_0, pixels_col_27_1, pixels_row_27_1, pixels_col_27_2, pixels_row_27_2, pixels_col_27_3, pixels_row_27_3, pixels_col_27_4, pixels_row_27_4, pixels_col_27_5, pixels_row_27_5, pixels_col_27_6, pixels_row_27_6, pixels_col_27_7, pixels_row_27_7, pixels_col_27_8, pixels_row_27_8, pixels_col_27_9, pixels_row_27_9, pixels_col_27_10, pixels_row_27_10, pixels_col_27_11, pixels_row_27_11, pixels_col_27_12, pixels_row_27_12, pixels_col_27_13, pixels_row_27_13, pixels_col_27_14, pixels_row_27_14, pixels_col_27_15, pixels_row_27_15, pixels_col_27_16, pixels_row_27_16, pixels_col_27_17, pixels_row_27_17, pixels_col_27_18, pixels_row_27_18, pixels_col_27_19, pixels_row_27_19, pixels_col_27_20, pixels_row_27_20, pixels_col_27_21, pixels_row_27_21, pixels_col_27_22, pixels_row_27_22, pixels_col_27_23, pixels_row_27_23, pixels_col_27_24, pixels_row_27_24, pixels_col_27_25, pixels_row_27_25, pixels_col_27_26, pixels_row_27_26, pixels_col_27_27, pixels_row_27_27, pixels_col_27_28, pixels_row_27_28, pixels_col_27_29, pixels_row_27_29, pixels_col_27_30, pixels_row_27_30, pixels_col_27_31, pixels_row_27_31, pixels_col_27_32, pixels_row_27_32, pixels_col_27_33, pixels_row_27_33, pixels_col_27_34, pixels_row_27_34, pixels_col_27_35, pixels_row_27_35, pixels_col_28_0, pixels_row_28_0, pixels_col_28_1, pixels_row_28_1, pixels_col_28_2, pixels_row_28_2, pixels_col_28_3, pixels_row_28_3, pixels_col_28_4, pixels_row_28_4, pixels_col_28_5, pixels_row_28_5, pixels_col_28_6, pixels_row_28_6, pixels_col_28_7, pixels_row_28_7, pixels_col_28_8, pixels_row_28_8, pixels_col_28_9, pixels_row_28_9, pixels_col_28_10, pixels_row_28_10, pixels_col_28_11, pixels_row_28_11, pixels_col_28_12, pixels_row_28_12, pixels_col_28_13, pixels_row_28_13, pixels_col_28_14, pixels_row_28_14, pixels_col_28_15, pixels_row_28_15, pixels_col_28_16, pixels_row_28_16, pixels_col_28_17, pixels_row_28_17, pixels_col_28_18, pixels_row_28_18, pixels_col_28_19, pixels_row_28_19, pixels_col_28_20, pixels_row_28_20, pixels_col_28_21, pixels_row_28_21, pixels_col_28_22, pixels_row_28_22, pixels_col_28_23, pixels_row_28_23, pixels_col_28_24, pixels_row_28_24, pixels_col_28_25, pixels_row_28_25, pixels_col_28_26, pixels_row_28_26, pixels_col_28_27, pixels_row_28_27, pixels_col_28_28, pixels_row_28_28, pixels_col_28_29, pixels_row_28_29, pixels_col_28_30, pixels_row_28_30, pixels_col_28_31, pixels_row_28_31, pixels_col_28_32, pixels_row_28_32, pixels_col_28_33, pixels_row_28_33, pixels_col_28_34, pixels_row_28_34, pixels_col_28_35, pixels_row_28_35, pixels_col_29_0, pixels_row_29_0, pixels_col_29_1, pixels_row_29_1, pixels_col_29_2, pixels_row_29_2, pixels_col_29_3, pixels_row_29_3, pixels_col_29_4, pixels_row_29_4, pixels_col_29_5, pixels_row_29_5, pixels_col_29_6, pixels_row_29_6, pixels_col_29_7, pixels_row_29_7, pixels_col_29_8, pixels_row_29_8, pixels_col_29_9, pixels_row_29_9, pixels_col_29_10, pixels_row_29_10, pixels_col_29_11, pixels_row_29_11, pixels_col_29_12, pixels_row_29_12, pixels_col_29_13, pixels_row_29_13, pixels_col_29_14, pixels_row_29_14, pixels_col_29_15, pixels_row_29_15, pixels_col_29_16, pixels_row_29_16, pixels_col_29_17, pixels_row_29_17, pixels_col_29_18, pixels_row_29_18, pixels_col_29_19, pixels_row_29_19, pixels_col_29_20, pixels_row_29_20, pixels_col_29_21, pixels_row_29_21, pixels_col_29_22, pixels_row_29_22, pixels_col_29_23, pixels_row_29_23, pixels_col_29_24, pixels_row_29_24, pixels_col_29_25, pixels_row_29_25, pixels_col_29_26, pixels_row_29_26, pixels_col_29_27, pixels_row_29_27, pixels_col_29_28, pixels_row_29_28, pixels_col_29_29, pixels_row_29_29, pixels_col_29_30, pixels_row_29_30, pixels_col_29_31, pixels_row_29_31, pixels_col_29_32, pixels_row_29_32, pixels_col_29_33, pixels_row_29_33, pixels_col_29_34, pixels_row_29_34, pixels_col_29_35, pixels_row_29_35, pixels_col_30_0, pixels_row_30_0, pixels_col_30_1, pixels_row_30_1, pixels_col_30_2, pixels_row_30_2, pixels_col_30_3, pixels_row_30_3, pixels_col_30_4, pixels_row_30_4, pixels_col_30_5, pixels_row_30_5, pixels_col_30_6, pixels_row_30_6, pixels_col_30_7, pixels_row_30_7, pixels_col_30_8, pixels_row_30_8, pixels_col_30_9, pixels_row_30_9, pixels_col_30_10, pixels_row_30_10, pixels_col_30_11, pixels_row_30_11, pixels_col_30_12, pixels_row_30_12, pixels_col_30_13, pixels_row_30_13, pixels_col_30_14, pixels_row_30_14, pixels_col_30_15, pixels_row_30_15, pixels_col_30_16, pixels_row_30_16, pixels_col_30_17, pixels_row_30_17, pixels_col_30_18, pixels_row_30_18, pixels_col_30_19, pixels_row_30_19, pixels_col_30_20, pixels_row_30_20, pixels_col_30_21, pixels_row_30_21, pixels_col_30_22, pixels_row_30_22, pixels_col_30_23, pixels_row_30_23, pixels_col_30_24, pixels_row_30_24, pixels_col_30_25, pixels_row_30_25, pixels_col_30_26, pixels_row_30_26, pixels_col_30_27, pixels_row_30_27, pixels_col_30_28, pixels_row_30_28, pixels_col_30_29, pixels_row_30_29, pixels_col_30_30, pixels_row_30_30, pixels_col_30_31, pixels_row_30_31, pixels_col_30_32, pixels_row_30_32, pixels_col_30_33, pixels_row_30_33, pixels_col_30_34, pixels_row_30_34, pixels_col_30_35, pixels_row_30_35, pixels_col_31_0, pixels_row_31_0, pixels_col_31_1, pixels_row_31_1, pixels_col_31_2, pixels_row_31_2, pixels_col_31_3, pixels_row_31_3, pixels_col_31_4, pixels_row_31_4, pixels_col_31_5, pixels_row_31_5, pixels_col_31_6, pixels_row_31_6, pixels_col_31_7, pixels_row_31_7, pixels_col_31_8, pixels_row_31_8, pixels_col_31_9, pixels_row_31_9, pixels_col_31_10, pixels_row_31_10, pixels_col_31_11, pixels_row_31_11, pixels_col_31_12, pixels_row_31_12, pixels_col_31_13, pixels_row_31_13, pixels_col_31_14, pixels_row_31_14, pixels_col_31_15, pixels_row_31_15, pixels_col_31_16, pixels_row_31_16, pixels_col_31_17, pixels_row_31_17, pixels_col_31_18, pixels_row_31_18, pixels_col_31_19, pixels_row_31_19, pixels_col_31_20, pixels_row_31_20, pixels_col_31_21, pixels_row_31_21, pixels_col_31_22, pixels_row_31_22, pixels_col_31_23, pixels_row_31_23, pixels_col_31_24, pixels_row_31_24, pixels_col_31_25, pixels_row_31_25, pixels_col_31_26, pixels_row_31_26, pixels_col_31_27, pixels_row_31_27, pixels_col_31_28, pixels_row_31_28, pixels_col_31_29, pixels_row_31_29, pixels_col_31_30, 
pixels_row_31_30, pixels_col_31_31, pixels_row_31_31, pixels_col_31_32, pixels_row_31_32, pixels_col_31_33, pixels_row_31_33, pixels_col_31_34, pixels_row_31_34, pixels_col_31_35, pixels_row_31_35, pixels_col_32_0, pixels_row_32_0, pixels_col_32_1, pixels_row_32_1, pixels_col_32_2, pixels_row_32_2, pixels_col_32_3, pixels_row_32_3, pixels_col_32_4, pixels_row_32_4, pixels_col_32_5, pixels_row_32_5, pixels_col_32_6, pixels_row_32_6, pixels_col_32_7, pixels_row_32_7, pixels_col_32_8, pixels_row_32_8, pixels_col_32_9, pixels_row_32_9, pixels_col_32_10, pixels_row_32_10, pixels_col_32_11, pixels_row_32_11, pixels_col_32_12, pixels_row_32_12, pixels_col_32_13, pixels_row_32_13, pixels_col_32_14, pixels_row_32_14, pixels_col_32_15, pixels_row_32_15, pixels_col_32_16, pixels_row_32_16, pixels_col_32_17, pixels_row_32_17, pixels_col_32_18, pixels_row_32_18, pixels_col_32_19, pixels_row_32_19, pixels_col_32_20, pixels_row_32_20, pixels_col_32_21, pixels_row_32_21, pixels_col_32_22, pixels_row_32_22, pixels_col_32_23, pixels_row_32_23, pixels_col_32_24, pixels_row_32_24, pixels_col_32_25, pixels_row_32_25, pixels_col_32_26, pixels_row_32_26, pixels_col_32_27, pixels_row_32_27, pixels_col_32_28, pixels_row_32_28, pixels_col_32_29, pixels_row_32_29, pixels_col_32_30, pixels_row_32_30, pixels_col_32_31, pixels_row_32_31, pixels_col_32_32, pixels_row_32_32, pixels_col_32_33, pixels_row_32_33, pixels_col_32_34, pixels_row_32_34, pixels_col_32_35, pixels_row_32_35, pixels_col_33_0, pixels_row_33_0, pixels_col_33_1, pixels_row_33_1, pixels_col_33_2, pixels_row_33_2, pixels_col_33_3, pixels_row_33_3, pixels_col_33_4, pixels_row_33_4, pixels_col_33_5, pixels_row_33_5, pixels_col_33_6, pixels_row_33_6, pixels_col_33_7, pixels_row_33_7, pixels_col_33_8, pixels_row_33_8, pixels_col_33_9, pixels_row_33_9, pixels_col_33_10, pixels_row_33_10, pixels_col_33_11, pixels_row_33_11, pixels_col_33_12, pixels_row_33_12, pixels_col_33_13, pixels_row_33_13, pixels_col_33_14, pixels_row_33_14, pixels_col_33_15, pixels_row_33_15, pixels_col_33_16, pixels_row_33_16, pixels_col_33_17, pixels_row_33_17, pixels_col_33_18, pixels_row_33_18, pixels_col_33_19, pixels_row_33_19, pixels_col_33_20, pixels_row_33_20, pixels_col_33_21, pixels_row_33_21, pixels_col_33_22, pixels_row_33_22, pixels_col_33_23, pixels_row_33_23, pixels_col_33_24, pixels_row_33_24, pixels_col_33_25, pixels_row_33_25, pixels_col_33_26, pixels_row_33_26, pixels_col_33_27, pixels_row_33_27, pixels_col_33_28, pixels_row_33_28, pixels_col_33_29, pixels_row_33_29, pixels_col_33_30, pixels_row_33_30, pixels_col_33_31, pixels_row_33_31, pixels_col_33_32, pixels_row_33_32, pixels_col_33_33, pixels_row_33_33, pixels_col_33_34, pixels_row_33_34, pixels_col_33_35, pixels_row_33_35, pixels_col_34_0, pixels_row_34_0, pixels_col_34_1, pixels_row_34_1, pixels_col_34_2, pixels_row_34_2, pixels_col_34_3, pixels_row_34_3, pixels_col_34_4, pixels_row_34_4, pixels_col_34_5, pixels_row_34_5, pixels_col_34_6, pixels_row_34_6, pixels_col_34_7, pixels_row_34_7, pixels_col_34_8, pixels_row_34_8, pixels_col_34_9, pixels_row_34_9, pixels_col_34_10, pixels_row_34_10, pixels_col_34_11, pixels_row_34_11, pixels_col_34_12, pixels_row_34_12, pixels_col_34_13, pixels_row_34_13, pixels_col_34_14, pixels_row_34_14, pixels_col_34_15, pixels_row_34_15, pixels_col_34_16, pixels_row_34_16, pixels_col_34_17, pixels_row_34_17, pixels_col_34_18, pixels_row_34_18, pixels_col_34_19, pixels_row_34_19, pixels_col_34_20, pixels_row_34_20, pixels_col_34_21, pixels_row_34_21, pixels_col_34_22, pixels_row_34_22, pixels_col_34_23, pixels_row_34_23, pixels_col_34_24, pixels_row_34_24, pixels_col_34_25, pixels_row_34_25, pixels_col_34_26, pixels_row_34_26, pixels_col_34_27, pixels_row_34_27, pixels_col_34_28, pixels_row_34_28, pixels_col_34_29, pixels_row_34_29, pixels_col_34_30, pixels_row_34_30, pixels_col_34_31, pixels_row_34_31, pixels_col_34_32, pixels_row_34_32, pixels_col_34_33, pixels_row_34_33, pixels_col_34_34, pixels_row_34_34, pixels_col_34_35, pixels_row_34_35, pixels_col_35_0, pixels_row_35_0, pixels_col_35_1, pixels_row_35_1, pixels_col_35_2, pixels_row_35_2, pixels_col_35_3, pixels_row_35_3, pixels_col_35_4, pixels_row_35_4, pixels_col_35_5, pixels_row_35_5, pixels_col_35_6, pixels_row_35_6, pixels_col_35_7, pixels_row_35_7, pixels_col_35_8, pixels_row_35_8, pixels_col_35_9, pixels_row_35_9, pixels_col_35_10, pixels_row_35_10, pixels_col_35_11, pixels_row_35_11, pixels_col_35_12, pixels_row_35_12, pixels_col_35_13, pixels_row_35_13, pixels_col_35_14, pixels_row_35_14, pixels_col_35_15, pixels_row_35_15, pixels_col_35_16, pixels_row_35_16, pixels_col_35_17, pixels_row_35_17, pixels_col_35_18, pixels_row_35_18, pixels_col_35_19, pixels_row_35_19, pixels_col_35_20, pixels_row_35_20, pixels_col_35_21, pixels_row_35_21, pixels_col_35_22, pixels_row_35_22, pixels_col_35_23, pixels_row_35_23, pixels_col_35_24, pixels_row_35_24, pixels_col_35_25, pixels_row_35_25, pixels_col_35_26, pixels_row_35_26, pixels_col_35_27, pixels_row_35_27, pixels_col_35_28, pixels_row_35_28, pixels_col_35_29, pixels_row_35_29, pixels_col_35_30, pixels_row_35_30, pixels_col_35_31, pixels_row_35_31, pixels_col_35_32, pixels_row_35_32, pixels_col_35_33, pixels_row_35_33, pixels_col_35_34, pixels_row_35_34, pixels_col_35_35, pixels_row_35_35;

assign pixels_col_0_0 = {data_out_cols[1*col_length-1 -: col_length]};
assign pixels_row_0_0 = {data_out_rows[1*col_length-1 -: col_length]};
assign pixels_col_0_1 = {data_out_cols[2*col_length-1 -: col_length]};
assign pixels_row_0_1 = {data_out_rows[2*col_length-1 -: col_length]};
assign pixels_col_0_2 = {data_out_cols[3*col_length-1 -: col_length]};
assign pixels_row_0_2 = {data_out_rows[3*col_length-1 -: col_length]};
assign pixels_col_0_3 = {data_out_cols[4*col_length-1 -: col_length]};
assign pixels_row_0_3 = {data_out_rows[4*col_length-1 -: col_length]};
assign pixels_col_0_4 = {data_out_cols[5*col_length-1 -: col_length]};
assign pixels_row_0_4 = {data_out_rows[5*col_length-1 -: col_length]};
assign pixels_col_0_5 = {data_out_cols[6*col_length-1 -: col_length]};
assign pixels_row_0_5 = {data_out_rows[6*col_length-1 -: col_length]};
assign pixels_col_0_6 = {data_out_cols[7*col_length-1 -: col_length]};
assign pixels_row_0_6 = {data_out_rows[7*col_length-1 -: col_length]};
assign pixels_col_0_7 = {data_out_cols[8*col_length-1 -: col_length]};
assign pixels_row_0_7 = {data_out_rows[8*col_length-1 -: col_length]};
assign pixels_col_0_8 = {data_out_cols[9*col_length-1 -: col_length]};
assign pixels_row_0_8 = {data_out_rows[9*col_length-1 -: col_length]};
assign pixels_col_0_9 = {data_out_cols[10*col_length-1 -: col_length]};
assign pixels_row_0_9 = {data_out_rows[10*col_length-1 -: col_length]};
assign pixels_col_0_10 = {data_out_cols[11*col_length-1 -: col_length]};
assign pixels_row_0_10 = {data_out_rows[11*col_length-1 -: col_length]};
assign pixels_col_0_11 = {data_out_cols[12*col_length-1 -: col_length]};
assign pixels_row_0_11 = {data_out_rows[12*col_length-1 -: col_length]};
assign pixels_col_0_12 = {data_out_cols[13*col_length-1 -: col_length]};
assign pixels_row_0_12 = {data_out_rows[13*col_length-1 -: col_length]};
assign pixels_col_0_13 = {data_out_cols[14*col_length-1 -: col_length]};
assign pixels_row_0_13 = {data_out_rows[14*col_length-1 -: col_length]};
assign pixels_col_0_14 = {data_out_cols[15*col_length-1 -: col_length]};
assign pixels_row_0_14 = {data_out_rows[15*col_length-1 -: col_length]};
assign pixels_col_0_15 = {data_out_cols[16*col_length-1 -: col_length]};
assign pixels_row_0_15 = {data_out_rows[16*col_length-1 -: col_length]};
assign pixels_col_0_16 = {data_out_cols[17*col_length-1 -: col_length]};
assign pixels_row_0_16 = {data_out_rows[17*col_length-1 -: col_length]};
assign pixels_col_0_17 = {data_out_cols[18*col_length-1 -: col_length]};
assign pixels_row_0_17 = {data_out_rows[18*col_length-1 -: col_length]};
assign pixels_col_0_18 = {data_out_cols[19*col_length-1 -: col_length]};
assign pixels_row_0_18 = {data_out_rows[19*col_length-1 -: col_length]};
assign pixels_col_0_19 = {data_out_cols[20*col_length-1 -: col_length]};
assign pixels_row_0_19 = {data_out_rows[20*col_length-1 -: col_length]};
assign pixels_col_0_20 = {data_out_cols[21*col_length-1 -: col_length]};
assign pixels_row_0_20 = {data_out_rows[21*col_length-1 -: col_length]};
assign pixels_col_0_21 = {data_out_cols[22*col_length-1 -: col_length]};
assign pixels_row_0_21 = {data_out_rows[22*col_length-1 -: col_length]};
assign pixels_col_0_22 = {data_out_cols[23*col_length-1 -: col_length]};
assign pixels_row_0_22 = {data_out_rows[23*col_length-1 -: col_length]};
assign pixels_col_0_23 = {data_out_cols[24*col_length-1 -: col_length]};
assign pixels_row_0_23 = {data_out_rows[24*col_length-1 -: col_length]};
assign pixels_col_0_24 = {data_out_cols[25*col_length-1 -: col_length]};
assign pixels_row_0_24 = {data_out_rows[25*col_length-1 -: col_length]};
assign pixels_col_0_25 = {data_out_cols[26*col_length-1 -: col_length]};
assign pixels_row_0_25 = {data_out_rows[26*col_length-1 -: col_length]};
assign pixels_col_0_26 = {data_out_cols[27*col_length-1 -: col_length]};
assign pixels_row_0_26 = {data_out_rows[27*col_length-1 -: col_length]};
assign pixels_col_0_27 = {data_out_cols[28*col_length-1 -: col_length]};
assign pixels_row_0_27 = {data_out_rows[28*col_length-1 -: col_length]};
assign pixels_col_0_28 = {data_out_cols[29*col_length-1 -: col_length]};
assign pixels_row_0_28 = {data_out_rows[29*col_length-1 -: col_length]};
assign pixels_col_0_29 = {data_out_cols[30*col_length-1 -: col_length]};
assign pixels_row_0_29 = {data_out_rows[30*col_length-1 -: col_length]};
assign pixels_col_0_30 = {data_out_cols[31*col_length-1 -: col_length]};
assign pixels_row_0_30 = {data_out_rows[31*col_length-1 -: col_length]};
assign pixels_col_0_31 = {data_out_cols[32*col_length-1 -: col_length]};
assign pixels_row_0_31 = {data_out_rows[32*col_length-1 -: col_length]};
assign pixels_col_0_32 = {data_out_cols[33*col_length-1 -: col_length]};
assign pixels_row_0_32 = {data_out_rows[33*col_length-1 -: col_length]};
assign pixels_col_0_33 = {data_out_cols[34*col_length-1 -: col_length]};
assign pixels_row_0_33 = {data_out_rows[34*col_length-1 -: col_length]};
assign pixels_col_0_34 = {data_out_cols[35*col_length-1 -: col_length]};
assign pixels_row_0_34 = {data_out_rows[35*col_length-1 -: col_length]};
assign pixels_col_0_35 = {data_out_cols[36*col_length-1 -: col_length]};
assign pixels_row_0_35 = {data_out_rows[36*col_length-1 -: col_length]};
assign pixels_col_1_0 = {data_out_cols[37*col_length-1 -: col_length]};
assign pixels_row_1_0 = {data_out_rows[37*col_length-1 -: col_length]};
assign pixels_col_1_1 = {data_out_cols[38*col_length-1 -: col_length]};
assign pixels_row_1_1 = {data_out_rows[38*col_length-1 -: col_length]};
assign pixels_col_1_2 = {data_out_cols[39*col_length-1 -: col_length]};
assign pixels_row_1_2 = {data_out_rows[39*col_length-1 -: col_length]};
assign pixels_col_1_3 = {data_out_cols[40*col_length-1 -: col_length]};
assign pixels_row_1_3 = {data_out_rows[40*col_length-1 -: col_length]};
assign pixels_col_1_4 = {data_out_cols[41*col_length-1 -: col_length]};
assign pixels_row_1_4 = {data_out_rows[41*col_length-1 -: col_length]};
assign pixels_col_1_5 = {data_out_cols[42*col_length-1 -: col_length]};
assign pixels_row_1_5 = {data_out_rows[42*col_length-1 -: col_length]};
assign pixels_col_1_6 = {data_out_cols[43*col_length-1 -: col_length]};
assign pixels_row_1_6 = {data_out_rows[43*col_length-1 -: col_length]};
assign pixels_col_1_7 = {data_out_cols[44*col_length-1 -: col_length]};
assign pixels_row_1_7 = {data_out_rows[44*col_length-1 -: col_length]};
assign pixels_col_1_8 = {data_out_cols[45*col_length-1 -: col_length]};
assign pixels_row_1_8 = {data_out_rows[45*col_length-1 -: col_length]};
assign pixels_col_1_9 = {data_out_cols[46*col_length-1 -: col_length]};
assign pixels_row_1_9 = {data_out_rows[46*col_length-1 -: col_length]};
assign pixels_col_1_10 = {data_out_cols[47*col_length-1 -: col_length]};
assign pixels_row_1_10 = {data_out_rows[47*col_length-1 -: col_length]};
assign pixels_col_1_11 = {data_out_cols[48*col_length-1 -: col_length]};
assign pixels_row_1_11 = {data_out_rows[48*col_length-1 -: col_length]};
assign pixels_col_1_12 = {data_out_cols[49*col_length-1 -: col_length]};
assign pixels_row_1_12 = {data_out_rows[49*col_length-1 -: col_length]};
assign pixels_col_1_13 = {data_out_cols[50*col_length-1 -: col_length]};
assign pixels_row_1_13 = {data_out_rows[50*col_length-1 -: col_length]};
assign pixels_col_1_14 = {data_out_cols[51*col_length-1 -: col_length]};
assign pixels_row_1_14 = {data_out_rows[51*col_length-1 -: col_length]};
assign pixels_col_1_15 = {data_out_cols[52*col_length-1 -: col_length]};
assign pixels_row_1_15 = {data_out_rows[52*col_length-1 -: col_length]};
assign pixels_col_1_16 = {data_out_cols[53*col_length-1 -: col_length]};
assign pixels_row_1_16 = {data_out_rows[53*col_length-1 -: col_length]};
assign pixels_col_1_17 = {data_out_cols[54*col_length-1 -: col_length]};
assign pixels_row_1_17 = {data_out_rows[54*col_length-1 -: col_length]};
assign pixels_col_1_18 = {data_out_cols[55*col_length-1 -: col_length]};
assign pixels_row_1_18 = {data_out_rows[55*col_length-1 -: col_length]};
assign pixels_col_1_19 = {data_out_cols[56*col_length-1 -: col_length]};
assign pixels_row_1_19 = {data_out_rows[56*col_length-1 -: col_length]};
assign pixels_col_1_20 = {data_out_cols[57*col_length-1 -: col_length]};
assign pixels_row_1_20 = {data_out_rows[57*col_length-1 -: col_length]};
assign pixels_col_1_21 = {data_out_cols[58*col_length-1 -: col_length]};
assign pixels_row_1_21 = {data_out_rows[58*col_length-1 -: col_length]};
assign pixels_col_1_22 = {data_out_cols[59*col_length-1 -: col_length]};
assign pixels_row_1_22 = {data_out_rows[59*col_length-1 -: col_length]};
assign pixels_col_1_23 = {data_out_cols[60*col_length-1 -: col_length]};
assign pixels_row_1_23 = {data_out_rows[60*col_length-1 -: col_length]};
assign pixels_col_1_24 = {data_out_cols[61*col_length-1 -: col_length]};
assign pixels_row_1_24 = {data_out_rows[61*col_length-1 -: col_length]};
assign pixels_col_1_25 = {data_out_cols[62*col_length-1 -: col_length]};
assign pixels_row_1_25 = {data_out_rows[62*col_length-1 -: col_length]};
assign pixels_col_1_26 = {data_out_cols[63*col_length-1 -: col_length]};
assign pixels_row_1_26 = {data_out_rows[63*col_length-1 -: col_length]};
assign pixels_col_1_27 = {data_out_cols[64*col_length-1 -: col_length]};
assign pixels_row_1_27 = {data_out_rows[64*col_length-1 -: col_length]};
assign pixels_col_1_28 = {data_out_cols[65*col_length-1 -: col_length]};
assign pixels_row_1_28 = {data_out_rows[65*col_length-1 -: col_length]};
assign pixels_col_1_29 = {data_out_cols[66*col_length-1 -: col_length]};
assign pixels_row_1_29 = {data_out_rows[66*col_length-1 -: col_length]};
assign pixels_col_1_30 = {data_out_cols[67*col_length-1 -: col_length]};
assign pixels_row_1_30 = {data_out_rows[67*col_length-1 -: col_length]};
assign pixels_col_1_31 = {data_out_cols[68*col_length-1 -: col_length]};
assign pixels_row_1_31 = {data_out_rows[68*col_length-1 -: col_length]};
assign pixels_col_1_32 = {data_out_cols[69*col_length-1 -: col_length]};
assign pixels_row_1_32 = {data_out_rows[69*col_length-1 -: col_length]};
assign pixels_col_1_33 = {data_out_cols[70*col_length-1 -: col_length]};
assign pixels_row_1_33 = {data_out_rows[70*col_length-1 -: col_length]};
assign pixels_col_1_34 = {data_out_cols[71*col_length-1 -: col_length]};
assign pixels_row_1_34 = {data_out_rows[71*col_length-1 -: col_length]};
assign pixels_col_1_35 = {data_out_cols[72*col_length-1 -: col_length]};
assign pixels_row_1_35 = {data_out_rows[72*col_length-1 -: col_length]};
assign pixels_col_2_0 = {data_out_cols[73*col_length-1 -: col_length]};
assign pixels_row_2_0 = {data_out_rows[73*col_length-1 -: col_length]};
assign pixels_col_2_1 = {data_out_cols[74*col_length-1 -: col_length]};
assign pixels_row_2_1 = {data_out_rows[74*col_length-1 -: col_length]};
assign pixels_col_2_2 = {data_out_cols[75*col_length-1 -: col_length]};
assign pixels_row_2_2 = {data_out_rows[75*col_length-1 -: col_length]};
assign pixels_col_2_3 = {data_out_cols[76*col_length-1 -: col_length]};
assign pixels_row_2_3 = {data_out_rows[76*col_length-1 -: col_length]};
assign pixels_col_2_4 = {data_out_cols[77*col_length-1 -: col_length]};
assign pixels_row_2_4 = {data_out_rows[77*col_length-1 -: col_length]};
assign pixels_col_2_5 = {data_out_cols[78*col_length-1 -: col_length]};
assign pixels_row_2_5 = {data_out_rows[78*col_length-1 -: col_length]};
assign pixels_col_2_6 = {data_out_cols[79*col_length-1 -: col_length]};
assign pixels_row_2_6 = {data_out_rows[79*col_length-1 -: col_length]};
assign pixels_col_2_7 = {data_out_cols[80*col_length-1 -: col_length]};
assign pixels_row_2_7 = {data_out_rows[80*col_length-1 -: col_length]};
assign pixels_col_2_8 = {data_out_cols[81*col_length-1 -: col_length]};
assign pixels_row_2_8 = {data_out_rows[81*col_length-1 -: col_length]};
assign pixels_col_2_9 = {data_out_cols[82*col_length-1 -: col_length]};
assign pixels_row_2_9 = {data_out_rows[82*col_length-1 -: col_length]};
assign pixels_col_2_10 = {data_out_cols[83*col_length-1 -: col_length]};
assign pixels_row_2_10 = {data_out_rows[83*col_length-1 -: col_length]};
assign pixels_col_2_11 = {data_out_cols[84*col_length-1 -: col_length]};
assign pixels_row_2_11 = {data_out_rows[84*col_length-1 -: col_length]};
assign pixels_col_2_12 = {data_out_cols[85*col_length-1 -: col_length]};
assign pixels_row_2_12 = {data_out_rows[85*col_length-1 -: col_length]};
assign pixels_col_2_13 = {data_out_cols[86*col_length-1 -: col_length]};
assign pixels_row_2_13 = {data_out_rows[86*col_length-1 -: col_length]};
assign pixels_col_2_14 = {data_out_cols[87*col_length-1 -: col_length]};
assign pixels_row_2_14 = {data_out_rows[87*col_length-1 -: col_length]};
assign pixels_col_2_15 = {data_out_cols[88*col_length-1 -: col_length]};
assign pixels_row_2_15 = {data_out_rows[88*col_length-1 -: col_length]};
assign pixels_col_2_16 = {data_out_cols[89*col_length-1 -: col_length]};
assign pixels_row_2_16 = {data_out_rows[89*col_length-1 -: col_length]};
assign pixels_col_2_17 = {data_out_cols[90*col_length-1 -: col_length]};
assign pixels_row_2_17 = {data_out_rows[90*col_length-1 -: col_length]};
assign pixels_col_2_18 = {data_out_cols[91*col_length-1 -: col_length]};
assign pixels_row_2_18 = {data_out_rows[91*col_length-1 -: col_length]};
assign pixels_col_2_19 = {data_out_cols[92*col_length-1 -: col_length]};
assign pixels_row_2_19 = {data_out_rows[92*col_length-1 -: col_length]};
assign pixels_col_2_20 = {data_out_cols[93*col_length-1 -: col_length]};
assign pixels_row_2_20 = {data_out_rows[93*col_length-1 -: col_length]};
assign pixels_col_2_21 = {data_out_cols[94*col_length-1 -: col_length]};
assign pixels_row_2_21 = {data_out_rows[94*col_length-1 -: col_length]};
assign pixels_col_2_22 = {data_out_cols[95*col_length-1 -: col_length]};
assign pixels_row_2_22 = {data_out_rows[95*col_length-1 -: col_length]};
assign pixels_col_2_23 = {data_out_cols[96*col_length-1 -: col_length]};
assign pixels_row_2_23 = {data_out_rows[96*col_length-1 -: col_length]};
assign pixels_col_2_24 = {data_out_cols[97*col_length-1 -: col_length]};
assign pixels_row_2_24 = {data_out_rows[97*col_length-1 -: col_length]};
assign pixels_col_2_25 = {data_out_cols[98*col_length-1 -: col_length]};
assign pixels_row_2_25 = {data_out_rows[98*col_length-1 -: col_length]};
assign pixels_col_2_26 = {data_out_cols[99*col_length-1 -: col_length]};
assign pixels_row_2_26 = {data_out_rows[99*col_length-1 -: col_length]};
assign pixels_col_2_27 = {data_out_cols[100*col_length-1 -: col_length]};
assign pixels_row_2_27 = {data_out_rows[100*col_length-1 -: col_length]};
assign pixels_col_2_28 = {data_out_cols[101*col_length-1 -: col_length]};
assign pixels_row_2_28 = {data_out_rows[101*col_length-1 -: col_length]};
assign pixels_col_2_29 = {data_out_cols[102*col_length-1 -: col_length]};
assign pixels_row_2_29 = {data_out_rows[102*col_length-1 -: col_length]};
assign pixels_col_2_30 = {data_out_cols[103*col_length-1 -: col_length]};
assign pixels_row_2_30 = {data_out_rows[103*col_length-1 -: col_length]};
assign pixels_col_2_31 = {data_out_cols[104*col_length-1 -: col_length]};
assign pixels_row_2_31 = {data_out_rows[104*col_length-1 -: col_length]};
assign pixels_col_2_32 = {data_out_cols[105*col_length-1 -: col_length]};
assign pixels_row_2_32 = {data_out_rows[105*col_length-1 -: col_length]};
assign pixels_col_2_33 = {data_out_cols[106*col_length-1 -: col_length]};
assign pixels_row_2_33 = {data_out_rows[106*col_length-1 -: col_length]};
assign pixels_col_2_34 = {data_out_cols[107*col_length-1 -: col_length]};
assign pixels_row_2_34 = {data_out_rows[107*col_length-1 -: col_length]};
assign pixels_col_2_35 = {data_out_cols[108*col_length-1 -: col_length]};
assign pixels_row_2_35 = {data_out_rows[108*col_length-1 -: col_length]};
assign pixels_col_3_0 = {data_out_cols[109*col_length-1 -: col_length]};
assign pixels_row_3_0 = {data_out_rows[109*col_length-1 -: col_length]};
assign pixels_col_3_1 = {data_out_cols[110*col_length-1 -: col_length]};
assign pixels_row_3_1 = {data_out_rows[110*col_length-1 -: col_length]};
assign pixels_col_3_2 = {data_out_cols[111*col_length-1 -: col_length]};
assign pixels_row_3_2 = {data_out_rows[111*col_length-1 -: col_length]};
assign pixels_col_3_3 = {data_out_cols[112*col_length-1 -: col_length]};
assign pixels_row_3_3 = {data_out_rows[112*col_length-1 -: col_length]};
assign pixels_col_3_4 = {data_out_cols[113*col_length-1 -: col_length]};
assign pixels_row_3_4 = {data_out_rows[113*col_length-1 -: col_length]};
assign pixels_col_3_5 = {data_out_cols[114*col_length-1 -: col_length]};
assign pixels_row_3_5 = {data_out_rows[114*col_length-1 -: col_length]};
assign pixels_col_3_6 = {data_out_cols[115*col_length-1 -: col_length]};
assign pixels_row_3_6 = {data_out_rows[115*col_length-1 -: col_length]};
assign pixels_col_3_7 = {data_out_cols[116*col_length-1 -: col_length]};
assign pixels_row_3_7 = {data_out_rows[116*col_length-1 -: col_length]};
assign pixels_col_3_8 = {data_out_cols[117*col_length-1 -: col_length]};
assign pixels_row_3_8 = {data_out_rows[117*col_length-1 -: col_length]};
assign pixels_col_3_9 = {data_out_cols[118*col_length-1 -: col_length]};
assign pixels_row_3_9 = {data_out_rows[118*col_length-1 -: col_length]};
assign pixels_col_3_10 = {data_out_cols[119*col_length-1 -: col_length]};
assign pixels_row_3_10 = {data_out_rows[119*col_length-1 -: col_length]};
assign pixels_col_3_11 = {data_out_cols[120*col_length-1 -: col_length]};
assign pixels_row_3_11 = {data_out_rows[120*col_length-1 -: col_length]};
assign pixels_col_3_12 = {data_out_cols[121*col_length-1 -: col_length]};
assign pixels_row_3_12 = {data_out_rows[121*col_length-1 -: col_length]};
assign pixels_col_3_13 = {data_out_cols[122*col_length-1 -: col_length]};
assign pixels_row_3_13 = {data_out_rows[122*col_length-1 -: col_length]};
assign pixels_col_3_14 = {data_out_cols[123*col_length-1 -: col_length]};
assign pixels_row_3_14 = {data_out_rows[123*col_length-1 -: col_length]};
assign pixels_col_3_15 = {data_out_cols[124*col_length-1 -: col_length]};
assign pixels_row_3_15 = {data_out_rows[124*col_length-1 -: col_length]};
assign pixels_col_3_16 = {data_out_cols[125*col_length-1 -: col_length]};
assign pixels_row_3_16 = {data_out_rows[125*col_length-1 -: col_length]};
assign pixels_col_3_17 = {data_out_cols[126*col_length-1 -: col_length]};
assign pixels_row_3_17 = {data_out_rows[126*col_length-1 -: col_length]};
assign pixels_col_3_18 = {data_out_cols[127*col_length-1 -: col_length]};
assign pixels_row_3_18 = {data_out_rows[127*col_length-1 -: col_length]};
assign pixels_col_3_19 = {data_out_cols[128*col_length-1 -: col_length]};
assign pixels_row_3_19 = {data_out_rows[128*col_length-1 -: col_length]};
assign pixels_col_3_20 = {data_out_cols[129*col_length-1 -: col_length]};
assign pixels_row_3_20 = {data_out_rows[129*col_length-1 -: col_length]};
assign pixels_col_3_21 = {data_out_cols[130*col_length-1 -: col_length]};
assign pixels_row_3_21 = {data_out_rows[130*col_length-1 -: col_length]};
assign pixels_col_3_22 = {data_out_cols[131*col_length-1 -: col_length]};
assign pixels_row_3_22 = {data_out_rows[131*col_length-1 -: col_length]};
assign pixels_col_3_23 = {data_out_cols[132*col_length-1 -: col_length]};
assign pixels_row_3_23 = {data_out_rows[132*col_length-1 -: col_length]};
assign pixels_col_3_24 = {data_out_cols[133*col_length-1 -: col_length]};
assign pixels_row_3_24 = {data_out_rows[133*col_length-1 -: col_length]};
assign pixels_col_3_25 = {data_out_cols[134*col_length-1 -: col_length]};
assign pixels_row_3_25 = {data_out_rows[134*col_length-1 -: col_length]};
assign pixels_col_3_26 = {data_out_cols[135*col_length-1 -: col_length]};
assign pixels_row_3_26 = {data_out_rows[135*col_length-1 -: col_length]};
assign pixels_col_3_27 = {data_out_cols[136*col_length-1 -: col_length]};
assign pixels_row_3_27 = {data_out_rows[136*col_length-1 -: col_length]};
assign pixels_col_3_28 = {data_out_cols[137*col_length-1 -: col_length]};
assign pixels_row_3_28 = {data_out_rows[137*col_length-1 -: col_length]};
assign pixels_col_3_29 = {data_out_cols[138*col_length-1 -: col_length]};
assign pixels_row_3_29 = {data_out_rows[138*col_length-1 -: col_length]};
assign pixels_col_3_30 = {data_out_cols[139*col_length-1 -: col_length]};
assign pixels_row_3_30 = {data_out_rows[139*col_length-1 -: col_length]};
assign pixels_col_3_31 = {data_out_cols[140*col_length-1 -: col_length]};
assign pixels_row_3_31 = {data_out_rows[140*col_length-1 -: col_length]};
assign pixels_col_3_32 = {data_out_cols[141*col_length-1 -: col_length]};
assign pixels_row_3_32 = {data_out_rows[141*col_length-1 -: col_length]};
assign pixels_col_3_33 = {data_out_cols[142*col_length-1 -: col_length]};
assign pixels_row_3_33 = {data_out_rows[142*col_length-1 -: col_length]};
assign pixels_col_3_34 = {data_out_cols[143*col_length-1 -: col_length]};
assign pixels_row_3_34 = {data_out_rows[143*col_length-1 -: col_length]};
assign pixels_col_3_35 = {data_out_cols[144*col_length-1 -: col_length]};
assign pixels_row_3_35 = {data_out_rows[144*col_length-1 -: col_length]};
assign pixels_col_4_0 = {data_out_cols[145*col_length-1 -: col_length]};
assign pixels_row_4_0 = {data_out_rows[145*col_length-1 -: col_length]};
assign pixels_col_4_1 = {data_out_cols[146*col_length-1 -: col_length]};
assign pixels_row_4_1 = {data_out_rows[146*col_length-1 -: col_length]};
assign pixels_col_4_2 = {data_out_cols[147*col_length-1 -: col_length]};
assign pixels_row_4_2 = {data_out_rows[147*col_length-1 -: col_length]};
assign pixels_col_4_3 = {data_out_cols[148*col_length-1 -: col_length]};
assign pixels_row_4_3 = {data_out_rows[148*col_length-1 -: col_length]};
assign pixels_col_4_4 = {data_out_cols[149*col_length-1 -: col_length]};
assign pixels_row_4_4 = {data_out_rows[149*col_length-1 -: col_length]};
assign pixels_col_4_5 = {data_out_cols[150*col_length-1 -: col_length]};
assign pixels_row_4_5 = {data_out_rows[150*col_length-1 -: col_length]};
assign pixels_col_4_6 = {data_out_cols[151*col_length-1 -: col_length]};
assign pixels_row_4_6 = {data_out_rows[151*col_length-1 -: col_length]};
assign pixels_col_4_7 = {data_out_cols[152*col_length-1 -: col_length]};
assign pixels_row_4_7 = {data_out_rows[152*col_length-1 -: col_length]};
assign pixels_col_4_8 = {data_out_cols[153*col_length-1 -: col_length]};
assign pixels_row_4_8 = {data_out_rows[153*col_length-1 -: col_length]};
assign pixels_col_4_9 = {data_out_cols[154*col_length-1 -: col_length]};
assign pixels_row_4_9 = {data_out_rows[154*col_length-1 -: col_length]};
assign pixels_col_4_10 = {data_out_cols[155*col_length-1 -: col_length]};
assign pixels_row_4_10 = {data_out_rows[155*col_length-1 -: col_length]};
assign pixels_col_4_11 = {data_out_cols[156*col_length-1 -: col_length]};
assign pixels_row_4_11 = {data_out_rows[156*col_length-1 -: col_length]};
assign pixels_col_4_12 = {data_out_cols[157*col_length-1 -: col_length]};
assign pixels_row_4_12 = {data_out_rows[157*col_length-1 -: col_length]};
assign pixels_col_4_13 = {data_out_cols[158*col_length-1 -: col_length]};
assign pixels_row_4_13 = {data_out_rows[158*col_length-1 -: col_length]};
assign pixels_col_4_14 = {data_out_cols[159*col_length-1 -: col_length]};
assign pixels_row_4_14 = {data_out_rows[159*col_length-1 -: col_length]};
assign pixels_col_4_15 = {data_out_cols[160*col_length-1 -: col_length]};
assign pixels_row_4_15 = {data_out_rows[160*col_length-1 -: col_length]};
assign pixels_col_4_16 = {data_out_cols[161*col_length-1 -: col_length]};
assign pixels_row_4_16 = {data_out_rows[161*col_length-1 -: col_length]};
assign pixels_col_4_17 = {data_out_cols[162*col_length-1 -: col_length]};
assign pixels_row_4_17 = {data_out_rows[162*col_length-1 -: col_length]};
assign pixels_col_4_18 = {data_out_cols[163*col_length-1 -: col_length]};
assign pixels_row_4_18 = {data_out_rows[163*col_length-1 -: col_length]};
assign pixels_col_4_19 = {data_out_cols[164*col_length-1 -: col_length]};
assign pixels_row_4_19 = {data_out_rows[164*col_length-1 -: col_length]};
assign pixels_col_4_20 = {data_out_cols[165*col_length-1 -: col_length]};
assign pixels_row_4_20 = {data_out_rows[165*col_length-1 -: col_length]};
assign pixels_col_4_21 = {data_out_cols[166*col_length-1 -: col_length]};
assign pixels_row_4_21 = {data_out_rows[166*col_length-1 -: col_length]};
assign pixels_col_4_22 = {data_out_cols[167*col_length-1 -: col_length]};
assign pixels_row_4_22 = {data_out_rows[167*col_length-1 -: col_length]};
assign pixels_col_4_23 = {data_out_cols[168*col_length-1 -: col_length]};
assign pixels_row_4_23 = {data_out_rows[168*col_length-1 -: col_length]};
assign pixels_col_4_24 = {data_out_cols[169*col_length-1 -: col_length]};
assign pixels_row_4_24 = {data_out_rows[169*col_length-1 -: col_length]};
assign pixels_col_4_25 = {data_out_cols[170*col_length-1 -: col_length]};
assign pixels_row_4_25 = {data_out_rows[170*col_length-1 -: col_length]};
assign pixels_col_4_26 = {data_out_cols[171*col_length-1 -: col_length]};
assign pixels_row_4_26 = {data_out_rows[171*col_length-1 -: col_length]};
assign pixels_col_4_27 = {data_out_cols[172*col_length-1 -: col_length]};
assign pixels_row_4_27 = {data_out_rows[172*col_length-1 -: col_length]};
assign pixels_col_4_28 = {data_out_cols[173*col_length-1 -: col_length]};
assign pixels_row_4_28 = {data_out_rows[173*col_length-1 -: col_length]};
assign pixels_col_4_29 = {data_out_cols[174*col_length-1 -: col_length]};
assign pixels_row_4_29 = {data_out_rows[174*col_length-1 -: col_length]};
assign pixels_col_4_30 = {data_out_cols[175*col_length-1 -: col_length]};
assign pixels_row_4_30 = {data_out_rows[175*col_length-1 -: col_length]};
assign pixels_col_4_31 = {data_out_cols[176*col_length-1 -: col_length]};
assign pixels_row_4_31 = {data_out_rows[176*col_length-1 -: col_length]};
assign pixels_col_4_32 = {data_out_cols[177*col_length-1 -: col_length]};
assign pixels_row_4_32 = {data_out_rows[177*col_length-1 -: col_length]};
assign pixels_col_4_33 = {data_out_cols[178*col_length-1 -: col_length]};
assign pixels_row_4_33 = {data_out_rows[178*col_length-1 -: col_length]};
assign pixels_col_4_34 = {data_out_cols[179*col_length-1 -: col_length]};
assign pixels_row_4_34 = {data_out_rows[179*col_length-1 -: col_length]};
assign pixels_col_4_35 = {data_out_cols[180*col_length-1 -: col_length]};
assign pixels_row_4_35 = {data_out_rows[180*col_length-1 -: col_length]};
assign pixels_col_5_0 = {data_out_cols[181*col_length-1 -: col_length]};
assign pixels_row_5_0 = {data_out_rows[181*col_length-1 -: col_length]};
assign pixels_col_5_1 = {data_out_cols[182*col_length-1 -: col_length]};
assign pixels_row_5_1 = {data_out_rows[182*col_length-1 -: col_length]};
assign pixels_col_5_2 = {data_out_cols[183*col_length-1 -: col_length]};
assign pixels_row_5_2 = {data_out_rows[183*col_length-1 -: col_length]};
assign pixels_col_5_3 = {data_out_cols[184*col_length-1 -: col_length]};
assign pixels_row_5_3 = {data_out_rows[184*col_length-1 -: col_length]};
assign pixels_col_5_4 = {data_out_cols[185*col_length-1 -: col_length]};
assign pixels_row_5_4 = {data_out_rows[185*col_length-1 -: col_length]};
assign pixels_col_5_5 = {data_out_cols[186*col_length-1 -: col_length]};
assign pixels_row_5_5 = {data_out_rows[186*col_length-1 -: col_length]};
assign pixels_col_5_6 = {data_out_cols[187*col_length-1 -: col_length]};
assign pixels_row_5_6 = {data_out_rows[187*col_length-1 -: col_length]};
assign pixels_col_5_7 = {data_out_cols[188*col_length-1 -: col_length]};
assign pixels_row_5_7 = {data_out_rows[188*col_length-1 -: col_length]};
assign pixels_col_5_8 = {data_out_cols[189*col_length-1 -: col_length]};
assign pixels_row_5_8 = {data_out_rows[189*col_length-1 -: col_length]};
assign pixels_col_5_9 = {data_out_cols[190*col_length-1 -: col_length]};
assign pixels_row_5_9 = {data_out_rows[190*col_length-1 -: col_length]};
assign pixels_col_5_10 = {data_out_cols[191*col_length-1 -: col_length]};
assign pixels_row_5_10 = {data_out_rows[191*col_length-1 -: col_length]};
assign pixels_col_5_11 = {data_out_cols[192*col_length-1 -: col_length]};
assign pixels_row_5_11 = {data_out_rows[192*col_length-1 -: col_length]};
assign pixels_col_5_12 = {data_out_cols[193*col_length-1 -: col_length]};
assign pixels_row_5_12 = {data_out_rows[193*col_length-1 -: col_length]};
assign pixels_col_5_13 = {data_out_cols[194*col_length-1 -: col_length]};
assign pixels_row_5_13 = {data_out_rows[194*col_length-1 -: col_length]};
assign pixels_col_5_14 = {data_out_cols[195*col_length-1 -: col_length]};
assign pixels_row_5_14 = {data_out_rows[195*col_length-1 -: col_length]};
assign pixels_col_5_15 = {data_out_cols[196*col_length-1 -: col_length]};
assign pixels_row_5_15 = {data_out_rows[196*col_length-1 -: col_length]};
assign pixels_col_5_16 = {data_out_cols[197*col_length-1 -: col_length]};
assign pixels_row_5_16 = {data_out_rows[197*col_length-1 -: col_length]};
assign pixels_col_5_17 = {data_out_cols[198*col_length-1 -: col_length]};
assign pixels_row_5_17 = {data_out_rows[198*col_length-1 -: col_length]};
assign pixels_col_5_18 = {data_out_cols[199*col_length-1 -: col_length]};
assign pixels_row_5_18 = {data_out_rows[199*col_length-1 -: col_length]};
assign pixels_col_5_19 = {data_out_cols[200*col_length-1 -: col_length]};
assign pixels_row_5_19 = {data_out_rows[200*col_length-1 -: col_length]};
assign pixels_col_5_20 = {data_out_cols[201*col_length-1 -: col_length]};
assign pixels_row_5_20 = {data_out_rows[201*col_length-1 -: col_length]};
assign pixels_col_5_21 = {data_out_cols[202*col_length-1 -: col_length]};
assign pixels_row_5_21 = {data_out_rows[202*col_length-1 -: col_length]};
assign pixels_col_5_22 = {data_out_cols[203*col_length-1 -: col_length]};
assign pixels_row_5_22 = {data_out_rows[203*col_length-1 -: col_length]};
assign pixels_col_5_23 = {data_out_cols[204*col_length-1 -: col_length]};
assign pixels_row_5_23 = {data_out_rows[204*col_length-1 -: col_length]};
assign pixels_col_5_24 = {data_out_cols[205*col_length-1 -: col_length]};
assign pixels_row_5_24 = {data_out_rows[205*col_length-1 -: col_length]};
assign pixels_col_5_25 = {data_out_cols[206*col_length-1 -: col_length]};
assign pixels_row_5_25 = {data_out_rows[206*col_length-1 -: col_length]};
assign pixels_col_5_26 = {data_out_cols[207*col_length-1 -: col_length]};
assign pixels_row_5_26 = {data_out_rows[207*col_length-1 -: col_length]};
assign pixels_col_5_27 = {data_out_cols[208*col_length-1 -: col_length]};
assign pixels_row_5_27 = {data_out_rows[208*col_length-1 -: col_length]};
assign pixels_col_5_28 = {data_out_cols[209*col_length-1 -: col_length]};
assign pixels_row_5_28 = {data_out_rows[209*col_length-1 -: col_length]};
assign pixels_col_5_29 = {data_out_cols[210*col_length-1 -: col_length]};
assign pixels_row_5_29 = {data_out_rows[210*col_length-1 -: col_length]};
assign pixels_col_5_30 = {data_out_cols[211*col_length-1 -: col_length]};
assign pixels_row_5_30 = {data_out_rows[211*col_length-1 -: col_length]};
assign pixels_col_5_31 = {data_out_cols[212*col_length-1 -: col_length]};
assign pixels_row_5_31 = {data_out_rows[212*col_length-1 -: col_length]};
assign pixels_col_5_32 = {data_out_cols[213*col_length-1 -: col_length]};
assign pixels_row_5_32 = {data_out_rows[213*col_length-1 -: col_length]};
assign pixels_col_5_33 = {data_out_cols[214*col_length-1 -: col_length]};
assign pixels_row_5_33 = {data_out_rows[214*col_length-1 -: col_length]};
assign pixels_col_5_34 = {data_out_cols[215*col_length-1 -: col_length]};
assign pixels_row_5_34 = {data_out_rows[215*col_length-1 -: col_length]};
assign pixels_col_5_35 = {data_out_cols[216*col_length-1 -: col_length]};
assign pixels_row_5_35 = {data_out_rows[216*col_length-1 -: col_length]};
assign pixels_col_6_0 = {data_out_cols[217*col_length-1 -: col_length]};
assign pixels_row_6_0 = {data_out_rows[217*col_length-1 -: col_length]};
assign pixels_col_6_1 = {data_out_cols[218*col_length-1 -: col_length]};
assign pixels_row_6_1 = {data_out_rows[218*col_length-1 -: col_length]};
assign pixels_col_6_2 = {data_out_cols[219*col_length-1 -: col_length]};
assign pixels_row_6_2 = {data_out_rows[219*col_length-1 -: col_length]};
assign pixels_col_6_3 = {data_out_cols[220*col_length-1 -: col_length]};
assign pixels_row_6_3 = {data_out_rows[220*col_length-1 -: col_length]};
assign pixels_col_6_4 = {data_out_cols[221*col_length-1 -: col_length]};
assign pixels_row_6_4 = {data_out_rows[221*col_length-1 -: col_length]};
assign pixels_col_6_5 = {data_out_cols[222*col_length-1 -: col_length]};
assign pixels_row_6_5 = {data_out_rows[222*col_length-1 -: col_length]};
assign pixels_col_6_6 = {data_out_cols[223*col_length-1 -: col_length]};
assign pixels_row_6_6 = {data_out_rows[223*col_length-1 -: col_length]};
assign pixels_col_6_7 = {data_out_cols[224*col_length-1 -: col_length]};
assign pixels_row_6_7 = {data_out_rows[224*col_length-1 -: col_length]};
assign pixels_col_6_8 = {data_out_cols[225*col_length-1 -: col_length]};
assign pixels_row_6_8 = {data_out_rows[225*col_length-1 -: col_length]};
assign pixels_col_6_9 = {data_out_cols[226*col_length-1 -: col_length]};
assign pixels_row_6_9 = {data_out_rows[226*col_length-1 -: col_length]};
assign pixels_col_6_10 = {data_out_cols[227*col_length-1 -: col_length]};
assign pixels_row_6_10 = {data_out_rows[227*col_length-1 -: col_length]};
assign pixels_col_6_11 = {data_out_cols[228*col_length-1 -: col_length]};
assign pixels_row_6_11 = {data_out_rows[228*col_length-1 -: col_length]};
assign pixels_col_6_12 = {data_out_cols[229*col_length-1 -: col_length]};
assign pixels_row_6_12 = {data_out_rows[229*col_length-1 -: col_length]};
assign pixels_col_6_13 = {data_out_cols[230*col_length-1 -: col_length]};
assign pixels_row_6_13 = {data_out_rows[230*col_length-1 -: col_length]};
assign pixels_col_6_14 = {data_out_cols[231*col_length-1 -: col_length]};
assign pixels_row_6_14 = {data_out_rows[231*col_length-1 -: col_length]};
assign pixels_col_6_15 = {data_out_cols[232*col_length-1 -: col_length]};
assign pixels_row_6_15 = {data_out_rows[232*col_length-1 -: col_length]};
assign pixels_col_6_16 = {data_out_cols[233*col_length-1 -: col_length]};
assign pixels_row_6_16 = {data_out_rows[233*col_length-1 -: col_length]};
assign pixels_col_6_17 = {data_out_cols[234*col_length-1 -: col_length]};
assign pixels_row_6_17 = {data_out_rows[234*col_length-1 -: col_length]};
assign pixels_col_6_18 = {data_out_cols[235*col_length-1 -: col_length]};
assign pixels_row_6_18 = {data_out_rows[235*col_length-1 -: col_length]};
assign pixels_col_6_19 = {data_out_cols[236*col_length-1 -: col_length]};
assign pixels_row_6_19 = {data_out_rows[236*col_length-1 -: col_length]};
assign pixels_col_6_20 = {data_out_cols[237*col_length-1 -: col_length]};
assign pixels_row_6_20 = {data_out_rows[237*col_length-1 -: col_length]};
assign pixels_col_6_21 = {data_out_cols[238*col_length-1 -: col_length]};
assign pixels_row_6_21 = {data_out_rows[238*col_length-1 -: col_length]};
assign pixels_col_6_22 = {data_out_cols[239*col_length-1 -: col_length]};
assign pixels_row_6_22 = {data_out_rows[239*col_length-1 -: col_length]};
assign pixels_col_6_23 = {data_out_cols[240*col_length-1 -: col_length]};
assign pixels_row_6_23 = {data_out_rows[240*col_length-1 -: col_length]};
assign pixels_col_6_24 = {data_out_cols[241*col_length-1 -: col_length]};
assign pixels_row_6_24 = {data_out_rows[241*col_length-1 -: col_length]};
assign pixels_col_6_25 = {data_out_cols[242*col_length-1 -: col_length]};
assign pixels_row_6_25 = {data_out_rows[242*col_length-1 -: col_length]};
assign pixels_col_6_26 = {data_out_cols[243*col_length-1 -: col_length]};
assign pixels_row_6_26 = {data_out_rows[243*col_length-1 -: col_length]};
assign pixels_col_6_27 = {data_out_cols[244*col_length-1 -: col_length]};
assign pixels_row_6_27 = {data_out_rows[244*col_length-1 -: col_length]};
assign pixels_col_6_28 = {data_out_cols[245*col_length-1 -: col_length]};
assign pixels_row_6_28 = {data_out_rows[245*col_length-1 -: col_length]};
assign pixels_col_6_29 = {data_out_cols[246*col_length-1 -: col_length]};
assign pixels_row_6_29 = {data_out_rows[246*col_length-1 -: col_length]};
assign pixels_col_6_30 = {data_out_cols[247*col_length-1 -: col_length]};
assign pixels_row_6_30 = {data_out_rows[247*col_length-1 -: col_length]};
assign pixels_col_6_31 = {data_out_cols[248*col_length-1 -: col_length]};
assign pixels_row_6_31 = {data_out_rows[248*col_length-1 -: col_length]};
assign pixels_col_6_32 = {data_out_cols[249*col_length-1 -: col_length]};
assign pixels_row_6_32 = {data_out_rows[249*col_length-1 -: col_length]};
assign pixels_col_6_33 = {data_out_cols[250*col_length-1 -: col_length]};
assign pixels_row_6_33 = {data_out_rows[250*col_length-1 -: col_length]};
assign pixels_col_6_34 = {data_out_cols[251*col_length-1 -: col_length]};
assign pixels_row_6_34 = {data_out_rows[251*col_length-1 -: col_length]};
assign pixels_col_6_35 = {data_out_cols[252*col_length-1 -: col_length]};
assign pixels_row_6_35 = {data_out_rows[252*col_length-1 -: col_length]};
assign pixels_col_7_0 = {data_out_cols[253*col_length-1 -: col_length]};
assign pixels_row_7_0 = {data_out_rows[253*col_length-1 -: col_length]};
assign pixels_col_7_1 = {data_out_cols[254*col_length-1 -: col_length]};
assign pixels_row_7_1 = {data_out_rows[254*col_length-1 -: col_length]};
assign pixels_col_7_2 = {data_out_cols[255*col_length-1 -: col_length]};
assign pixels_row_7_2 = {data_out_rows[255*col_length-1 -: col_length]};
assign pixels_col_7_3 = {data_out_cols[256*col_length-1 -: col_length]};
assign pixels_row_7_3 = {data_out_rows[256*col_length-1 -: col_length]};
assign pixels_col_7_4 = {data_out_cols[257*col_length-1 -: col_length]};
assign pixels_row_7_4 = {data_out_rows[257*col_length-1 -: col_length]};
assign pixels_col_7_5 = {data_out_cols[258*col_length-1 -: col_length]};
assign pixels_row_7_5 = {data_out_rows[258*col_length-1 -: col_length]};
assign pixels_col_7_6 = {data_out_cols[259*col_length-1 -: col_length]};
assign pixels_row_7_6 = {data_out_rows[259*col_length-1 -: col_length]};
assign pixels_col_7_7 = {data_out_cols[260*col_length-1 -: col_length]};
assign pixels_row_7_7 = {data_out_rows[260*col_length-1 -: col_length]};
assign pixels_col_7_8 = {data_out_cols[261*col_length-1 -: col_length]};
assign pixels_row_7_8 = {data_out_rows[261*col_length-1 -: col_length]};
assign pixels_col_7_9 = {data_out_cols[262*col_length-1 -: col_length]};
assign pixels_row_7_9 = {data_out_rows[262*col_length-1 -: col_length]};
assign pixels_col_7_10 = {data_out_cols[263*col_length-1 -: col_length]};
assign pixels_row_7_10 = {data_out_rows[263*col_length-1 -: col_length]};
assign pixels_col_7_11 = {data_out_cols[264*col_length-1 -: col_length]};
assign pixels_row_7_11 = {data_out_rows[264*col_length-1 -: col_length]};
assign pixels_col_7_12 = {data_out_cols[265*col_length-1 -: col_length]};
assign pixels_row_7_12 = {data_out_rows[265*col_length-1 -: col_length]};
assign pixels_col_7_13 = {data_out_cols[266*col_length-1 -: col_length]};
assign pixels_row_7_13 = {data_out_rows[266*col_length-1 -: col_length]};
assign pixels_col_7_14 = {data_out_cols[267*col_length-1 -: col_length]};
assign pixels_row_7_14 = {data_out_rows[267*col_length-1 -: col_length]};
assign pixels_col_7_15 = {data_out_cols[268*col_length-1 -: col_length]};
assign pixels_row_7_15 = {data_out_rows[268*col_length-1 -: col_length]};
assign pixels_col_7_16 = {data_out_cols[269*col_length-1 -: col_length]};
assign pixels_row_7_16 = {data_out_rows[269*col_length-1 -: col_length]};
assign pixels_col_7_17 = {data_out_cols[270*col_length-1 -: col_length]};
assign pixels_row_7_17 = {data_out_rows[270*col_length-1 -: col_length]};
assign pixels_col_7_18 = {data_out_cols[271*col_length-1 -: col_length]};
assign pixels_row_7_18 = {data_out_rows[271*col_length-1 -: col_length]};
assign pixels_col_7_19 = {data_out_cols[272*col_length-1 -: col_length]};
assign pixels_row_7_19 = {data_out_rows[272*col_length-1 -: col_length]};
assign pixels_col_7_20 = {data_out_cols[273*col_length-1 -: col_length]};
assign pixels_row_7_20 = {data_out_rows[273*col_length-1 -: col_length]};
assign pixels_col_7_21 = {data_out_cols[274*col_length-1 -: col_length]};
assign pixels_row_7_21 = {data_out_rows[274*col_length-1 -: col_length]};
assign pixels_col_7_22 = {data_out_cols[275*col_length-1 -: col_length]};
assign pixels_row_7_22 = {data_out_rows[275*col_length-1 -: col_length]};
assign pixels_col_7_23 = {data_out_cols[276*col_length-1 -: col_length]};
assign pixels_row_7_23 = {data_out_rows[276*col_length-1 -: col_length]};
assign pixels_col_7_24 = {data_out_cols[277*col_length-1 -: col_length]};
assign pixels_row_7_24 = {data_out_rows[277*col_length-1 -: col_length]};
assign pixels_col_7_25 = {data_out_cols[278*col_length-1 -: col_length]};
assign pixels_row_7_25 = {data_out_rows[278*col_length-1 -: col_length]};
assign pixels_col_7_26 = {data_out_cols[279*col_length-1 -: col_length]};
assign pixels_row_7_26 = {data_out_rows[279*col_length-1 -: col_length]};
assign pixels_col_7_27 = {data_out_cols[280*col_length-1 -: col_length]};
assign pixels_row_7_27 = {data_out_rows[280*col_length-1 -: col_length]};
assign pixels_col_7_28 = {data_out_cols[281*col_length-1 -: col_length]};
assign pixels_row_7_28 = {data_out_rows[281*col_length-1 -: col_length]};
assign pixels_col_7_29 = {data_out_cols[282*col_length-1 -: col_length]};
assign pixels_row_7_29 = {data_out_rows[282*col_length-1 -: col_length]};
assign pixels_col_7_30 = {data_out_cols[283*col_length-1 -: col_length]};
assign pixels_row_7_30 = {data_out_rows[283*col_length-1 -: col_length]};
assign pixels_col_7_31 = {data_out_cols[284*col_length-1 -: col_length]};
assign pixels_row_7_31 = {data_out_rows[284*col_length-1 -: col_length]};
assign pixels_col_7_32 = {data_out_cols[285*col_length-1 -: col_length]};
assign pixels_row_7_32 = {data_out_rows[285*col_length-1 -: col_length]};
assign pixels_col_7_33 = {data_out_cols[286*col_length-1 -: col_length]};
assign pixels_row_7_33 = {data_out_rows[286*col_length-1 -: col_length]};
assign pixels_col_7_34 = {data_out_cols[287*col_length-1 -: col_length]};
assign pixels_row_7_34 = {data_out_rows[287*col_length-1 -: col_length]};
assign pixels_col_7_35 = {data_out_cols[288*col_length-1 -: col_length]};
assign pixels_row_7_35 = {data_out_rows[288*col_length-1 -: col_length]};
assign pixels_col_8_0 = {data_out_cols[289*col_length-1 -: col_length]};
assign pixels_row_8_0 = {data_out_rows[289*col_length-1 -: col_length]};
assign pixels_col_8_1 = {data_out_cols[290*col_length-1 -: col_length]};
assign pixels_row_8_1 = {data_out_rows[290*col_length-1 -: col_length]};
assign pixels_col_8_2 = {data_out_cols[291*col_length-1 -: col_length]};
assign pixels_row_8_2 = {data_out_rows[291*col_length-1 -: col_length]};
assign pixels_col_8_3 = {data_out_cols[292*col_length-1 -: col_length]};
assign pixels_row_8_3 = {data_out_rows[292*col_length-1 -: col_length]};
assign pixels_col_8_4 = {data_out_cols[293*col_length-1 -: col_length]};
assign pixels_row_8_4 = {data_out_rows[293*col_length-1 -: col_length]};
assign pixels_col_8_5 = {data_out_cols[294*col_length-1 -: col_length]};
assign pixels_row_8_5 = {data_out_rows[294*col_length-1 -: col_length]};
assign pixels_col_8_6 = {data_out_cols[295*col_length-1 -: col_length]};
assign pixels_row_8_6 = {data_out_rows[295*col_length-1 -: col_length]};
assign pixels_col_8_7 = {data_out_cols[296*col_length-1 -: col_length]};
assign pixels_row_8_7 = {data_out_rows[296*col_length-1 -: col_length]};
assign pixels_col_8_8 = {data_out_cols[297*col_length-1 -: col_length]};
assign pixels_row_8_8 = {data_out_rows[297*col_length-1 -: col_length]};
assign pixels_col_8_9 = {data_out_cols[298*col_length-1 -: col_length]};
assign pixels_row_8_9 = {data_out_rows[298*col_length-1 -: col_length]};
assign pixels_col_8_10 = {data_out_cols[299*col_length-1 -: col_length]};
assign pixels_row_8_10 = {data_out_rows[299*col_length-1 -: col_length]};
assign pixels_col_8_11 = {data_out_cols[300*col_length-1 -: col_length]};
assign pixels_row_8_11 = {data_out_rows[300*col_length-1 -: col_length]};
assign pixels_col_8_12 = {data_out_cols[301*col_length-1 -: col_length]};
assign pixels_row_8_12 = {data_out_rows[301*col_length-1 -: col_length]};
assign pixels_col_8_13 = {data_out_cols[302*col_length-1 -: col_length]};
assign pixels_row_8_13 = {data_out_rows[302*col_length-1 -: col_length]};
assign pixels_col_8_14 = {data_out_cols[303*col_length-1 -: col_length]};
assign pixels_row_8_14 = {data_out_rows[303*col_length-1 -: col_length]};
assign pixels_col_8_15 = {data_out_cols[304*col_length-1 -: col_length]};
assign pixels_row_8_15 = {data_out_rows[304*col_length-1 -: col_length]};
assign pixels_col_8_16 = {data_out_cols[305*col_length-1 -: col_length]};
assign pixels_row_8_16 = {data_out_rows[305*col_length-1 -: col_length]};
assign pixels_col_8_17 = {data_out_cols[306*col_length-1 -: col_length]};
assign pixels_row_8_17 = {data_out_rows[306*col_length-1 -: col_length]};
assign pixels_col_8_18 = {data_out_cols[307*col_length-1 -: col_length]};
assign pixels_row_8_18 = {data_out_rows[307*col_length-1 -: col_length]};
assign pixels_col_8_19 = {data_out_cols[308*col_length-1 -: col_length]};
assign pixels_row_8_19 = {data_out_rows[308*col_length-1 -: col_length]};
assign pixels_col_8_20 = {data_out_cols[309*col_length-1 -: col_length]};
assign pixels_row_8_20 = {data_out_rows[309*col_length-1 -: col_length]};
assign pixels_col_8_21 = {data_out_cols[310*col_length-1 -: col_length]};
assign pixels_row_8_21 = {data_out_rows[310*col_length-1 -: col_length]};
assign pixels_col_8_22 = {data_out_cols[311*col_length-1 -: col_length]};
assign pixels_row_8_22 = {data_out_rows[311*col_length-1 -: col_length]};
assign pixels_col_8_23 = {data_out_cols[312*col_length-1 -: col_length]};
assign pixels_row_8_23 = {data_out_rows[312*col_length-1 -: col_length]};
assign pixels_col_8_24 = {data_out_cols[313*col_length-1 -: col_length]};
assign pixels_row_8_24 = {data_out_rows[313*col_length-1 -: col_length]};
assign pixels_col_8_25 = {data_out_cols[314*col_length-1 -: col_length]};
assign pixels_row_8_25 = {data_out_rows[314*col_length-1 -: col_length]};
assign pixels_col_8_26 = {data_out_cols[315*col_length-1 -: col_length]};
assign pixels_row_8_26 = {data_out_rows[315*col_length-1 -: col_length]};
assign pixels_col_8_27 = {data_out_cols[316*col_length-1 -: col_length]};
assign pixels_row_8_27 = {data_out_rows[316*col_length-1 -: col_length]};
assign pixels_col_8_28 = {data_out_cols[317*col_length-1 -: col_length]};
assign pixels_row_8_28 = {data_out_rows[317*col_length-1 -: col_length]};
assign pixels_col_8_29 = {data_out_cols[318*col_length-1 -: col_length]};
assign pixels_row_8_29 = {data_out_rows[318*col_length-1 -: col_length]};
assign pixels_col_8_30 = {data_out_cols[319*col_length-1 -: col_length]};
assign pixels_row_8_30 = {data_out_rows[319*col_length-1 -: col_length]};
assign pixels_col_8_31 = {data_out_cols[320*col_length-1 -: col_length]};
assign pixels_row_8_31 = {data_out_rows[320*col_length-1 -: col_length]};
assign pixels_col_8_32 = {data_out_cols[321*col_length-1 -: col_length]};
assign pixels_row_8_32 = {data_out_rows[321*col_length-1 -: col_length]};
assign pixels_col_8_33 = {data_out_cols[322*col_length-1 -: col_length]};
assign pixels_row_8_33 = {data_out_rows[322*col_length-1 -: col_length]};
assign pixels_col_8_34 = {data_out_cols[323*col_length-1 -: col_length]};
assign pixels_row_8_34 = {data_out_rows[323*col_length-1 -: col_length]};
assign pixels_col_8_35 = {data_out_cols[324*col_length-1 -: col_length]};
assign pixels_row_8_35 = {data_out_rows[324*col_length-1 -: col_length]};
assign pixels_col_9_0 = {data_out_cols[325*col_length-1 -: col_length]};
assign pixels_row_9_0 = {data_out_rows[325*col_length-1 -: col_length]};
assign pixels_col_9_1 = {data_out_cols[326*col_length-1 -: col_length]};
assign pixels_row_9_1 = {data_out_rows[326*col_length-1 -: col_length]};
assign pixels_col_9_2 = {data_out_cols[327*col_length-1 -: col_length]};
assign pixels_row_9_2 = {data_out_rows[327*col_length-1 -: col_length]};
assign pixels_col_9_3 = {data_out_cols[328*col_length-1 -: col_length]};
assign pixels_row_9_3 = {data_out_rows[328*col_length-1 -: col_length]};
assign pixels_col_9_4 = {data_out_cols[329*col_length-1 -: col_length]};
assign pixels_row_9_4 = {data_out_rows[329*col_length-1 -: col_length]};
assign pixels_col_9_5 = {data_out_cols[330*col_length-1 -: col_length]};
assign pixels_row_9_5 = {data_out_rows[330*col_length-1 -: col_length]};
assign pixels_col_9_6 = {data_out_cols[331*col_length-1 -: col_length]};
assign pixels_row_9_6 = {data_out_rows[331*col_length-1 -: col_length]};
assign pixels_col_9_7 = {data_out_cols[332*col_length-1 -: col_length]};
assign pixels_row_9_7 = {data_out_rows[332*col_length-1 -: col_length]};
assign pixels_col_9_8 = {data_out_cols[333*col_length-1 -: col_length]};
assign pixels_row_9_8 = {data_out_rows[333*col_length-1 -: col_length]};
assign pixels_col_9_9 = {data_out_cols[334*col_length-1 -: col_length]};
assign pixels_row_9_9 = {data_out_rows[334*col_length-1 -: col_length]};
assign pixels_col_9_10 = {data_out_cols[335*col_length-1 -: col_length]};
assign pixels_row_9_10 = {data_out_rows[335*col_length-1 -: col_length]};
assign pixels_col_9_11 = {data_out_cols[336*col_length-1 -: col_length]};
assign pixels_row_9_11 = {data_out_rows[336*col_length-1 -: col_length]};
assign pixels_col_9_12 = {data_out_cols[337*col_length-1 -: col_length]};
assign pixels_row_9_12 = {data_out_rows[337*col_length-1 -: col_length]};
assign pixels_col_9_13 = {data_out_cols[338*col_length-1 -: col_length]};
assign pixels_row_9_13 = {data_out_rows[338*col_length-1 -: col_length]};
assign pixels_col_9_14 = {data_out_cols[339*col_length-1 -: col_length]};
assign pixels_row_9_14 = {data_out_rows[339*col_length-1 -: col_length]};
assign pixels_col_9_15 = {data_out_cols[340*col_length-1 -: col_length]};
assign pixels_row_9_15 = {data_out_rows[340*col_length-1 -: col_length]};
assign pixels_col_9_16 = {data_out_cols[341*col_length-1 -: col_length]};
assign pixels_row_9_16 = {data_out_rows[341*col_length-1 -: col_length]};
assign pixels_col_9_17 = {data_out_cols[342*col_length-1 -: col_length]};
assign pixels_row_9_17 = {data_out_rows[342*col_length-1 -: col_length]};
assign pixels_col_9_18 = {data_out_cols[343*col_length-1 -: col_length]};
assign pixels_row_9_18 = {data_out_rows[343*col_length-1 -: col_length]};
assign pixels_col_9_19 = {data_out_cols[344*col_length-1 -: col_length]};
assign pixels_row_9_19 = {data_out_rows[344*col_length-1 -: col_length]};
assign pixels_col_9_20 = {data_out_cols[345*col_length-1 -: col_length]};
assign pixels_row_9_20 = {data_out_rows[345*col_length-1 -: col_length]};
assign pixels_col_9_21 = {data_out_cols[346*col_length-1 -: col_length]};
assign pixels_row_9_21 = {data_out_rows[346*col_length-1 -: col_length]};
assign pixels_col_9_22 = {data_out_cols[347*col_length-1 -: col_length]};
assign pixels_row_9_22 = {data_out_rows[347*col_length-1 -: col_length]};
assign pixels_col_9_23 = {data_out_cols[348*col_length-1 -: col_length]};
assign pixels_row_9_23 = {data_out_rows[348*col_length-1 -: col_length]};
assign pixels_col_9_24 = {data_out_cols[349*col_length-1 -: col_length]};
assign pixels_row_9_24 = {data_out_rows[349*col_length-1 -: col_length]};
assign pixels_col_9_25 = {data_out_cols[350*col_length-1 -: col_length]};
assign pixels_row_9_25 = {data_out_rows[350*col_length-1 -: col_length]};
assign pixels_col_9_26 = {data_out_cols[351*col_length-1 -: col_length]};
assign pixels_row_9_26 = {data_out_rows[351*col_length-1 -: col_length]};
assign pixels_col_9_27 = {data_out_cols[352*col_length-1 -: col_length]};
assign pixels_row_9_27 = {data_out_rows[352*col_length-1 -: col_length]};
assign pixels_col_9_28 = {data_out_cols[353*col_length-1 -: col_length]};
assign pixels_row_9_28 = {data_out_rows[353*col_length-1 -: col_length]};
assign pixels_col_9_29 = {data_out_cols[354*col_length-1 -: col_length]};
assign pixels_row_9_29 = {data_out_rows[354*col_length-1 -: col_length]};
assign pixels_col_9_30 = {data_out_cols[355*col_length-1 -: col_length]};
assign pixels_row_9_30 = {data_out_rows[355*col_length-1 -: col_length]};
assign pixels_col_9_31 = {data_out_cols[356*col_length-1 -: col_length]};
assign pixels_row_9_31 = {data_out_rows[356*col_length-1 -: col_length]};
assign pixels_col_9_32 = {data_out_cols[357*col_length-1 -: col_length]};
assign pixels_row_9_32 = {data_out_rows[357*col_length-1 -: col_length]};
assign pixels_col_9_33 = {data_out_cols[358*col_length-1 -: col_length]};
assign pixels_row_9_33 = {data_out_rows[358*col_length-1 -: col_length]};
assign pixels_col_9_34 = {data_out_cols[359*col_length-1 -: col_length]};
assign pixels_row_9_34 = {data_out_rows[359*col_length-1 -: col_length]};
assign pixels_col_9_35 = {data_out_cols[360*col_length-1 -: col_length]};
assign pixels_row_9_35 = {data_out_rows[360*col_length-1 -: col_length]};
assign pixels_col_10_0 = {data_out_cols[361*col_length-1 -: col_length]};
assign pixels_row_10_0 = {data_out_rows[361*col_length-1 -: col_length]};
assign pixels_col_10_1 = {data_out_cols[362*col_length-1 -: col_length]};
assign pixels_row_10_1 = {data_out_rows[362*col_length-1 -: col_length]};
assign pixels_col_10_2 = {data_out_cols[363*col_length-1 -: col_length]};
assign pixels_row_10_2 = {data_out_rows[363*col_length-1 -: col_length]};
assign pixels_col_10_3 = {data_out_cols[364*col_length-1 -: col_length]};
assign pixels_row_10_3 = {data_out_rows[364*col_length-1 -: col_length]};
assign pixels_col_10_4 = {data_out_cols[365*col_length-1 -: col_length]};
assign pixels_row_10_4 = {data_out_rows[365*col_length-1 -: col_length]};
assign pixels_col_10_5 = {data_out_cols[366*col_length-1 -: col_length]};
assign pixels_row_10_5 = {data_out_rows[366*col_length-1 -: col_length]};
assign pixels_col_10_6 = {data_out_cols[367*col_length-1 -: col_length]};
assign pixels_row_10_6 = {data_out_rows[367*col_length-1 -: col_length]};
assign pixels_col_10_7 = {data_out_cols[368*col_length-1 -: col_length]};
assign pixels_row_10_7 = {data_out_rows[368*col_length-1 -: col_length]};
assign pixels_col_10_8 = {data_out_cols[369*col_length-1 -: col_length]};
assign pixels_row_10_8 = {data_out_rows[369*col_length-1 -: col_length]};
assign pixels_col_10_9 = {data_out_cols[370*col_length-1 -: col_length]};
assign pixels_row_10_9 = {data_out_rows[370*col_length-1 -: col_length]};
assign pixels_col_10_10 = {data_out_cols[371*col_length-1 -: col_length]};
assign pixels_row_10_10 = {data_out_rows[371*col_length-1 -: col_length]};
assign pixels_col_10_11 = {data_out_cols[372*col_length-1 -: col_length]};
assign pixels_row_10_11 = {data_out_rows[372*col_length-1 -: col_length]};
assign pixels_col_10_12 = {data_out_cols[373*col_length-1 -: col_length]};
assign pixels_row_10_12 = {data_out_rows[373*col_length-1 -: col_length]};
assign pixels_col_10_13 = {data_out_cols[374*col_length-1 -: col_length]};
assign pixels_row_10_13 = {data_out_rows[374*col_length-1 -: col_length]};
assign pixels_col_10_14 = {data_out_cols[375*col_length-1 -: col_length]};
assign pixels_row_10_14 = {data_out_rows[375*col_length-1 -: col_length]};
assign pixels_col_10_15 = {data_out_cols[376*col_length-1 -: col_length]};
assign pixels_row_10_15 = {data_out_rows[376*col_length-1 -: col_length]};
assign pixels_col_10_16 = {data_out_cols[377*col_length-1 -: col_length]};
assign pixels_row_10_16 = {data_out_rows[377*col_length-1 -: col_length]};
assign pixels_col_10_17 = {data_out_cols[378*col_length-1 -: col_length]};
assign pixels_row_10_17 = {data_out_rows[378*col_length-1 -: col_length]};
assign pixels_col_10_18 = {data_out_cols[379*col_length-1 -: col_length]};
assign pixels_row_10_18 = {data_out_rows[379*col_length-1 -: col_length]};
assign pixels_col_10_19 = {data_out_cols[380*col_length-1 -: col_length]};
assign pixels_row_10_19 = {data_out_rows[380*col_length-1 -: col_length]};
assign pixels_col_10_20 = {data_out_cols[381*col_length-1 -: col_length]};
assign pixels_row_10_20 = {data_out_rows[381*col_length-1 -: col_length]};
assign pixels_col_10_21 = {data_out_cols[382*col_length-1 -: col_length]};
assign pixels_row_10_21 = {data_out_rows[382*col_length-1 -: col_length]};
assign pixels_col_10_22 = {data_out_cols[383*col_length-1 -: col_length]};
assign pixels_row_10_22 = {data_out_rows[383*col_length-1 -: col_length]};
assign pixels_col_10_23 = {data_out_cols[384*col_length-1 -: col_length]};
assign pixels_row_10_23 = {data_out_rows[384*col_length-1 -: col_length]};
assign pixels_col_10_24 = {data_out_cols[385*col_length-1 -: col_length]};
assign pixels_row_10_24 = {data_out_rows[385*col_length-1 -: col_length]};
assign pixels_col_10_25 = {data_out_cols[386*col_length-1 -: col_length]};
assign pixels_row_10_25 = {data_out_rows[386*col_length-1 -: col_length]};
assign pixels_col_10_26 = {data_out_cols[387*col_length-1 -: col_length]};
assign pixels_row_10_26 = {data_out_rows[387*col_length-1 -: col_length]};
assign pixels_col_10_27 = {data_out_cols[388*col_length-1 -: col_length]};
assign pixels_row_10_27 = {data_out_rows[388*col_length-1 -: col_length]};
assign pixels_col_10_28 = {data_out_cols[389*col_length-1 -: col_length]};
assign pixels_row_10_28 = {data_out_rows[389*col_length-1 -: col_length]};
assign pixels_col_10_29 = {data_out_cols[390*col_length-1 -: col_length]};
assign pixels_row_10_29 = {data_out_rows[390*col_length-1 -: col_length]};
assign pixels_col_10_30 = {data_out_cols[391*col_length-1 -: col_length]};
assign pixels_row_10_30 = {data_out_rows[391*col_length-1 -: col_length]};
assign pixels_col_10_31 = {data_out_cols[392*col_length-1 -: col_length]};
assign pixels_row_10_31 = {data_out_rows[392*col_length-1 -: col_length]};
assign pixels_col_10_32 = {data_out_cols[393*col_length-1 -: col_length]};
assign pixels_row_10_32 = {data_out_rows[393*col_length-1 -: col_length]};
assign pixels_col_10_33 = {data_out_cols[394*col_length-1 -: col_length]};
assign pixels_row_10_33 = {data_out_rows[394*col_length-1 -: col_length]};
assign pixels_col_10_34 = {data_out_cols[395*col_length-1 -: col_length]};
assign pixels_row_10_34 = {data_out_rows[395*col_length-1 -: col_length]};
assign pixels_col_10_35 = {data_out_cols[396*col_length-1 -: col_length]};
assign pixels_row_10_35 = {data_out_rows[396*col_length-1 -: col_length]};
assign pixels_col_11_0 = {data_out_cols[397*col_length-1 -: col_length]};
assign pixels_row_11_0 = {data_out_rows[397*col_length-1 -: col_length]};
assign pixels_col_11_1 = {data_out_cols[398*col_length-1 -: col_length]};
assign pixels_row_11_1 = {data_out_rows[398*col_length-1 -: col_length]};
assign pixels_col_11_2 = {data_out_cols[399*col_length-1 -: col_length]};
assign pixels_row_11_2 = {data_out_rows[399*col_length-1 -: col_length]};
assign pixels_col_11_3 = {data_out_cols[400*col_length-1 -: col_length]};
assign pixels_row_11_3 = {data_out_rows[400*col_length-1 -: col_length]};
assign pixels_col_11_4 = {data_out_cols[401*col_length-1 -: col_length]};
assign pixels_row_11_4 = {data_out_rows[401*col_length-1 -: col_length]};
assign pixels_col_11_5 = {data_out_cols[402*col_length-1 -: col_length]};
assign pixels_row_11_5 = {data_out_rows[402*col_length-1 -: col_length]};
assign pixels_col_11_6 = {data_out_cols[403*col_length-1 -: col_length]};
assign pixels_row_11_6 = {data_out_rows[403*col_length-1 -: col_length]};
assign pixels_col_11_7 = {data_out_cols[404*col_length-1 -: col_length]};
assign pixels_row_11_7 = {data_out_rows[404*col_length-1 -: col_length]};
assign pixels_col_11_8 = {data_out_cols[405*col_length-1 -: col_length]};
assign pixels_row_11_8 = {data_out_rows[405*col_length-1 -: col_length]};
assign pixels_col_11_9 = {data_out_cols[406*col_length-1 -: col_length]};
assign pixels_row_11_9 = {data_out_rows[406*col_length-1 -: col_length]};
assign pixels_col_11_10 = {data_out_cols[407*col_length-1 -: col_length]};
assign pixels_row_11_10 = {data_out_rows[407*col_length-1 -: col_length]};
assign pixels_col_11_11 = {data_out_cols[408*col_length-1 -: col_length]};
assign pixels_row_11_11 = {data_out_rows[408*col_length-1 -: col_length]};
assign pixels_col_11_12 = {data_out_cols[409*col_length-1 -: col_length]};
assign pixels_row_11_12 = {data_out_rows[409*col_length-1 -: col_length]};
assign pixels_col_11_13 = {data_out_cols[410*col_length-1 -: col_length]};
assign pixels_row_11_13 = {data_out_rows[410*col_length-1 -: col_length]};
assign pixels_col_11_14 = {data_out_cols[411*col_length-1 -: col_length]};
assign pixels_row_11_14 = {data_out_rows[411*col_length-1 -: col_length]};
assign pixels_col_11_15 = {data_out_cols[412*col_length-1 -: col_length]};
assign pixels_row_11_15 = {data_out_rows[412*col_length-1 -: col_length]};
assign pixels_col_11_16 = {data_out_cols[413*col_length-1 -: col_length]};
assign pixels_row_11_16 = {data_out_rows[413*col_length-1 -: col_length]};
assign pixels_col_11_17 = {data_out_cols[414*col_length-1 -: col_length]};
assign pixels_row_11_17 = {data_out_rows[414*col_length-1 -: col_length]};
assign pixels_col_11_18 = {data_out_cols[415*col_length-1 -: col_length]};
assign pixels_row_11_18 = {data_out_rows[415*col_length-1 -: col_length]};
assign pixels_col_11_19 = {data_out_cols[416*col_length-1 -: col_length]};
assign pixels_row_11_19 = {data_out_rows[416*col_length-1 -: col_length]};
assign pixels_col_11_20 = {data_out_cols[417*col_length-1 -: col_length]};
assign pixels_row_11_20 = {data_out_rows[417*col_length-1 -: col_length]};
assign pixels_col_11_21 = {data_out_cols[418*col_length-1 -: col_length]};
assign pixels_row_11_21 = {data_out_rows[418*col_length-1 -: col_length]};
assign pixels_col_11_22 = {data_out_cols[419*col_length-1 -: col_length]};
assign pixels_row_11_22 = {data_out_rows[419*col_length-1 -: col_length]};
assign pixels_col_11_23 = {data_out_cols[420*col_length-1 -: col_length]};
assign pixels_row_11_23 = {data_out_rows[420*col_length-1 -: col_length]};
assign pixels_col_11_24 = {data_out_cols[421*col_length-1 -: col_length]};
assign pixels_row_11_24 = {data_out_rows[421*col_length-1 -: col_length]};
assign pixels_col_11_25 = {data_out_cols[422*col_length-1 -: col_length]};
assign pixels_row_11_25 = {data_out_rows[422*col_length-1 -: col_length]};
assign pixels_col_11_26 = {data_out_cols[423*col_length-1 -: col_length]};
assign pixels_row_11_26 = {data_out_rows[423*col_length-1 -: col_length]};
assign pixels_col_11_27 = {data_out_cols[424*col_length-1 -: col_length]};
assign pixels_row_11_27 = {data_out_rows[424*col_length-1 -: col_length]};
assign pixels_col_11_28 = {data_out_cols[425*col_length-1 -: col_length]};
assign pixels_row_11_28 = {data_out_rows[425*col_length-1 -: col_length]};
assign pixels_col_11_29 = {data_out_cols[426*col_length-1 -: col_length]};
assign pixels_row_11_29 = {data_out_rows[426*col_length-1 -: col_length]};
assign pixels_col_11_30 = {data_out_cols[427*col_length-1 -: col_length]};
assign pixels_row_11_30 = {data_out_rows[427*col_length-1 -: col_length]};
assign pixels_col_11_31 = {data_out_cols[428*col_length-1 -: col_length]};
assign pixels_row_11_31 = {data_out_rows[428*col_length-1 -: col_length]};
assign pixels_col_11_32 = {data_out_cols[429*col_length-1 -: col_length]};
assign pixels_row_11_32 = {data_out_rows[429*col_length-1 -: col_length]};
assign pixels_col_11_33 = {data_out_cols[430*col_length-1 -: col_length]};
assign pixels_row_11_33 = {data_out_rows[430*col_length-1 -: col_length]};
assign pixels_col_11_34 = {data_out_cols[431*col_length-1 -: col_length]};
assign pixels_row_11_34 = {data_out_rows[431*col_length-1 -: col_length]};
assign pixels_col_11_35 = {data_out_cols[432*col_length-1 -: col_length]};
assign pixels_row_11_35 = {data_out_rows[432*col_length-1 -: col_length]};
assign pixels_col_12_0 = {data_out_cols[433*col_length-1 -: col_length]};
assign pixels_row_12_0 = {data_out_rows[433*col_length-1 -: col_length]};
assign pixels_col_12_1 = {data_out_cols[434*col_length-1 -: col_length]};
assign pixels_row_12_1 = {data_out_rows[434*col_length-1 -: col_length]};
assign pixels_col_12_2 = {data_out_cols[435*col_length-1 -: col_length]};
assign pixels_row_12_2 = {data_out_rows[435*col_length-1 -: col_length]};
assign pixels_col_12_3 = {data_out_cols[436*col_length-1 -: col_length]};
assign pixels_row_12_3 = {data_out_rows[436*col_length-1 -: col_length]};
assign pixels_col_12_4 = {data_out_cols[437*col_length-1 -: col_length]};
assign pixels_row_12_4 = {data_out_rows[437*col_length-1 -: col_length]};
assign pixels_col_12_5 = {data_out_cols[438*col_length-1 -: col_length]};
assign pixels_row_12_5 = {data_out_rows[438*col_length-1 -: col_length]};
assign pixels_col_12_6 = {data_out_cols[439*col_length-1 -: col_length]};
assign pixels_row_12_6 = {data_out_rows[439*col_length-1 -: col_length]};
assign pixels_col_12_7 = {data_out_cols[440*col_length-1 -: col_length]};
assign pixels_row_12_7 = {data_out_rows[440*col_length-1 -: col_length]};
assign pixels_col_12_8 = {data_out_cols[441*col_length-1 -: col_length]};
assign pixels_row_12_8 = {data_out_rows[441*col_length-1 -: col_length]};
assign pixels_col_12_9 = {data_out_cols[442*col_length-1 -: col_length]};
assign pixels_row_12_9 = {data_out_rows[442*col_length-1 -: col_length]};
assign pixels_col_12_10 = {data_out_cols[443*col_length-1 -: col_length]};
assign pixels_row_12_10 = {data_out_rows[443*col_length-1 -: col_length]};
assign pixels_col_12_11 = {data_out_cols[444*col_length-1 -: col_length]};
assign pixels_row_12_11 = {data_out_rows[444*col_length-1 -: col_length]};
assign pixels_col_12_12 = {data_out_cols[445*col_length-1 -: col_length]};
assign pixels_row_12_12 = {data_out_rows[445*col_length-1 -: col_length]};
assign pixels_col_12_13 = {data_out_cols[446*col_length-1 -: col_length]};
assign pixels_row_12_13 = {data_out_rows[446*col_length-1 -: col_length]};
assign pixels_col_12_14 = {data_out_cols[447*col_length-1 -: col_length]};
assign pixels_row_12_14 = {data_out_rows[447*col_length-1 -: col_length]};
assign pixels_col_12_15 = {data_out_cols[448*col_length-1 -: col_length]};
assign pixels_row_12_15 = {data_out_rows[448*col_length-1 -: col_length]};
assign pixels_col_12_16 = {data_out_cols[449*col_length-1 -: col_length]};
assign pixels_row_12_16 = {data_out_rows[449*col_length-1 -: col_length]};
assign pixels_col_12_17 = {data_out_cols[450*col_length-1 -: col_length]};
assign pixels_row_12_17 = {data_out_rows[450*col_length-1 -: col_length]};
assign pixels_col_12_18 = {data_out_cols[451*col_length-1 -: col_length]};
assign pixels_row_12_18 = {data_out_rows[451*col_length-1 -: col_length]};
assign pixels_col_12_19 = {data_out_cols[452*col_length-1 -: col_length]};
assign pixels_row_12_19 = {data_out_rows[452*col_length-1 -: col_length]};
assign pixels_col_12_20 = {data_out_cols[453*col_length-1 -: col_length]};
assign pixels_row_12_20 = {data_out_rows[453*col_length-1 -: col_length]};
assign pixels_col_12_21 = {data_out_cols[454*col_length-1 -: col_length]};
assign pixels_row_12_21 = {data_out_rows[454*col_length-1 -: col_length]};
assign pixels_col_12_22 = {data_out_cols[455*col_length-1 -: col_length]};
assign pixels_row_12_22 = {data_out_rows[455*col_length-1 -: col_length]};
assign pixels_col_12_23 = {data_out_cols[456*col_length-1 -: col_length]};
assign pixels_row_12_23 = {data_out_rows[456*col_length-1 -: col_length]};
assign pixels_col_12_24 = {data_out_cols[457*col_length-1 -: col_length]};
assign pixels_row_12_24 = {data_out_rows[457*col_length-1 -: col_length]};
assign pixels_col_12_25 = {data_out_cols[458*col_length-1 -: col_length]};
assign pixels_row_12_25 = {data_out_rows[458*col_length-1 -: col_length]};
assign pixels_col_12_26 = {data_out_cols[459*col_length-1 -: col_length]};
assign pixels_row_12_26 = {data_out_rows[459*col_length-1 -: col_length]};
assign pixels_col_12_27 = {data_out_cols[460*col_length-1 -: col_length]};
assign pixels_row_12_27 = {data_out_rows[460*col_length-1 -: col_length]};
assign pixels_col_12_28 = {data_out_cols[461*col_length-1 -: col_length]};
assign pixels_row_12_28 = {data_out_rows[461*col_length-1 -: col_length]};
assign pixels_col_12_29 = {data_out_cols[462*col_length-1 -: col_length]};
assign pixels_row_12_29 = {data_out_rows[462*col_length-1 -: col_length]};
assign pixels_col_12_30 = {data_out_cols[463*col_length-1 -: col_length]};
assign pixels_row_12_30 = {data_out_rows[463*col_length-1 -: col_length]};
assign pixels_col_12_31 = {data_out_cols[464*col_length-1 -: col_length]};
assign pixels_row_12_31 = {data_out_rows[464*col_length-1 -: col_length]};
assign pixels_col_12_32 = {data_out_cols[465*col_length-1 -: col_length]};
assign pixels_row_12_32 = {data_out_rows[465*col_length-1 -: col_length]};
assign pixels_col_12_33 = {data_out_cols[466*col_length-1 -: col_length]};
assign pixels_row_12_33 = {data_out_rows[466*col_length-1 -: col_length]};
assign pixels_col_12_34 = {data_out_cols[467*col_length-1 -: col_length]};
assign pixels_row_12_34 = {data_out_rows[467*col_length-1 -: col_length]};
assign pixels_col_12_35 = {data_out_cols[468*col_length-1 -: col_length]};
assign pixels_row_12_35 = {data_out_rows[468*col_length-1 -: col_length]};
assign pixels_col_13_0 = {data_out_cols[469*col_length-1 -: col_length]};
assign pixels_row_13_0 = {data_out_rows[469*col_length-1 -: col_length]};
assign pixels_col_13_1 = {data_out_cols[470*col_length-1 -: col_length]};
assign pixels_row_13_1 = {data_out_rows[470*col_length-1 -: col_length]};
assign pixels_col_13_2 = {data_out_cols[471*col_length-1 -: col_length]};
assign pixels_row_13_2 = {data_out_rows[471*col_length-1 -: col_length]};
assign pixels_col_13_3 = {data_out_cols[472*col_length-1 -: col_length]};
assign pixels_row_13_3 = {data_out_rows[472*col_length-1 -: col_length]};
assign pixels_col_13_4 = {data_out_cols[473*col_length-1 -: col_length]};
assign pixels_row_13_4 = {data_out_rows[473*col_length-1 -: col_length]};
assign pixels_col_13_5 = {data_out_cols[474*col_length-1 -: col_length]};
assign pixels_row_13_5 = {data_out_rows[474*col_length-1 -: col_length]};
assign pixels_col_13_6 = {data_out_cols[475*col_length-1 -: col_length]};
assign pixels_row_13_6 = {data_out_rows[475*col_length-1 -: col_length]};
assign pixels_col_13_7 = {data_out_cols[476*col_length-1 -: col_length]};
assign pixels_row_13_7 = {data_out_rows[476*col_length-1 -: col_length]};
assign pixels_col_13_8 = {data_out_cols[477*col_length-1 -: col_length]};
assign pixels_row_13_8 = {data_out_rows[477*col_length-1 -: col_length]};
assign pixels_col_13_9 = {data_out_cols[478*col_length-1 -: col_length]};
assign pixels_row_13_9 = {data_out_rows[478*col_length-1 -: col_length]};
assign pixels_col_13_10 = {data_out_cols[479*col_length-1 -: col_length]};
assign pixels_row_13_10 = {data_out_rows[479*col_length-1 -: col_length]};
assign pixels_col_13_11 = {data_out_cols[480*col_length-1 -: col_length]};
assign pixels_row_13_11 = {data_out_rows[480*col_length-1 -: col_length]};
assign pixels_col_13_12 = {data_out_cols[481*col_length-1 -: col_length]};
assign pixels_row_13_12 = {data_out_rows[481*col_length-1 -: col_length]};
assign pixels_col_13_13 = {data_out_cols[482*col_length-1 -: col_length]};
assign pixels_row_13_13 = {data_out_rows[482*col_length-1 -: col_length]};
assign pixels_col_13_14 = {data_out_cols[483*col_length-1 -: col_length]};
assign pixels_row_13_14 = {data_out_rows[483*col_length-1 -: col_length]};
assign pixels_col_13_15 = {data_out_cols[484*col_length-1 -: col_length]};
assign pixels_row_13_15 = {data_out_rows[484*col_length-1 -: col_length]};
assign pixels_col_13_16 = {data_out_cols[485*col_length-1 -: col_length]};
assign pixels_row_13_16 = {data_out_rows[485*col_length-1 -: col_length]};
assign pixels_col_13_17 = {data_out_cols[486*col_length-1 -: col_length]};
assign pixels_row_13_17 = {data_out_rows[486*col_length-1 -: col_length]};
assign pixels_col_13_18 = {data_out_cols[487*col_length-1 -: col_length]};
assign pixels_row_13_18 = {data_out_rows[487*col_length-1 -: col_length]};
assign pixels_col_13_19 = {data_out_cols[488*col_length-1 -: col_length]};
assign pixels_row_13_19 = {data_out_rows[488*col_length-1 -: col_length]};
assign pixels_col_13_20 = {data_out_cols[489*col_length-1 -: col_length]};
assign pixels_row_13_20 = {data_out_rows[489*col_length-1 -: col_length]};
assign pixels_col_13_21 = {data_out_cols[490*col_length-1 -: col_length]};
assign pixels_row_13_21 = {data_out_rows[490*col_length-1 -: col_length]};
assign pixels_col_13_22 = {data_out_cols[491*col_length-1 -: col_length]};
assign pixels_row_13_22 = {data_out_rows[491*col_length-1 -: col_length]};
assign pixels_col_13_23 = {data_out_cols[492*col_length-1 -: col_length]};
assign pixels_row_13_23 = {data_out_rows[492*col_length-1 -: col_length]};
assign pixels_col_13_24 = {data_out_cols[493*col_length-1 -: col_length]};
assign pixels_row_13_24 = {data_out_rows[493*col_length-1 -: col_length]};
assign pixels_col_13_25 = {data_out_cols[494*col_length-1 -: col_length]};
assign pixels_row_13_25 = {data_out_rows[494*col_length-1 -: col_length]};
assign pixels_col_13_26 = {data_out_cols[495*col_length-1 -: col_length]};
assign pixels_row_13_26 = {data_out_rows[495*col_length-1 -: col_length]};
assign pixels_col_13_27 = {data_out_cols[496*col_length-1 -: col_length]};
assign pixels_row_13_27 = {data_out_rows[496*col_length-1 -: col_length]};
assign pixels_col_13_28 = {data_out_cols[497*col_length-1 -: col_length]};
assign pixels_row_13_28 = {data_out_rows[497*col_length-1 -: col_length]};
assign pixels_col_13_29 = {data_out_cols[498*col_length-1 -: col_length]};
assign pixels_row_13_29 = {data_out_rows[498*col_length-1 -: col_length]};
assign pixels_col_13_30 = {data_out_cols[499*col_length-1 -: col_length]};
assign pixels_row_13_30 = {data_out_rows[499*col_length-1 -: col_length]};
assign pixels_col_13_31 = {data_out_cols[500*col_length-1 -: col_length]};
assign pixels_row_13_31 = {data_out_rows[500*col_length-1 -: col_length]};
assign pixels_col_13_32 = {data_out_cols[501*col_length-1 -: col_length]};
assign pixels_row_13_32 = {data_out_rows[501*col_length-1 -: col_length]};
assign pixels_col_13_33 = {data_out_cols[502*col_length-1 -: col_length]};
assign pixels_row_13_33 = {data_out_rows[502*col_length-1 -: col_length]};
assign pixels_col_13_34 = {data_out_cols[503*col_length-1 -: col_length]};
assign pixels_row_13_34 = {data_out_rows[503*col_length-1 -: col_length]};
assign pixels_col_13_35 = {data_out_cols[504*col_length-1 -: col_length]};
assign pixels_row_13_35 = {data_out_rows[504*col_length-1 -: col_length]};
assign pixels_col_14_0 = {data_out_cols[505*col_length-1 -: col_length]};
assign pixels_row_14_0 = {data_out_rows[505*col_length-1 -: col_length]};
assign pixels_col_14_1 = {data_out_cols[506*col_length-1 -: col_length]};
assign pixels_row_14_1 = {data_out_rows[506*col_length-1 -: col_length]};
assign pixels_col_14_2 = {data_out_cols[507*col_length-1 -: col_length]};
assign pixels_row_14_2 = {data_out_rows[507*col_length-1 -: col_length]};
assign pixels_col_14_3 = {data_out_cols[508*col_length-1 -: col_length]};
assign pixels_row_14_3 = {data_out_rows[508*col_length-1 -: col_length]};
assign pixels_col_14_4 = {data_out_cols[509*col_length-1 -: col_length]};
assign pixels_row_14_4 = {data_out_rows[509*col_length-1 -: col_length]};
assign pixels_col_14_5 = {data_out_cols[510*col_length-1 -: col_length]};
assign pixels_row_14_5 = {data_out_rows[510*col_length-1 -: col_length]};
assign pixels_col_14_6 = {data_out_cols[511*col_length-1 -: col_length]};
assign pixels_row_14_6 = {data_out_rows[511*col_length-1 -: col_length]};
assign pixels_col_14_7 = {data_out_cols[512*col_length-1 -: col_length]};
assign pixels_row_14_7 = {data_out_rows[512*col_length-1 -: col_length]};
assign pixels_col_14_8 = {data_out_cols[513*col_length-1 -: col_length]};
assign pixels_row_14_8 = {data_out_rows[513*col_length-1 -: col_length]};
assign pixels_col_14_9 = {data_out_cols[514*col_length-1 -: col_length]};
assign pixels_row_14_9 = {data_out_rows[514*col_length-1 -: col_length]};
assign pixels_col_14_10 = {data_out_cols[515*col_length-1 -: col_length]};
assign pixels_row_14_10 = {data_out_rows[515*col_length-1 -: col_length]};
assign pixels_col_14_11 = {data_out_cols[516*col_length-1 -: col_length]};
assign pixels_row_14_11 = {data_out_rows[516*col_length-1 -: col_length]};
assign pixels_col_14_12 = {data_out_cols[517*col_length-1 -: col_length]};
assign pixels_row_14_12 = {data_out_rows[517*col_length-1 -: col_length]};
assign pixels_col_14_13 = {data_out_cols[518*col_length-1 -: col_length]};
assign pixels_row_14_13 = {data_out_rows[518*col_length-1 -: col_length]};
assign pixels_col_14_14 = {data_out_cols[519*col_length-1 -: col_length]};
assign pixels_row_14_14 = {data_out_rows[519*col_length-1 -: col_length]};
assign pixels_col_14_15 = {data_out_cols[520*col_length-1 -: col_length]};
assign pixels_row_14_15 = {data_out_rows[520*col_length-1 -: col_length]};
assign pixels_col_14_16 = {data_out_cols[521*col_length-1 -: col_length]};
assign pixels_row_14_16 = {data_out_rows[521*col_length-1 -: col_length]};
assign pixels_col_14_17 = {data_out_cols[522*col_length-1 -: col_length]};
assign pixels_row_14_17 = {data_out_rows[522*col_length-1 -: col_length]};
assign pixels_col_14_18 = {data_out_cols[523*col_length-1 -: col_length]};
assign pixels_row_14_18 = {data_out_rows[523*col_length-1 -: col_length]};
assign pixels_col_14_19 = {data_out_cols[524*col_length-1 -: col_length]};
assign pixels_row_14_19 = {data_out_rows[524*col_length-1 -: col_length]};
assign pixels_col_14_20 = {data_out_cols[525*col_length-1 -: col_length]};
assign pixels_row_14_20 = {data_out_rows[525*col_length-1 -: col_length]};
assign pixels_col_14_21 = {data_out_cols[526*col_length-1 -: col_length]};
assign pixels_row_14_21 = {data_out_rows[526*col_length-1 -: col_length]};
assign pixels_col_14_22 = {data_out_cols[527*col_length-1 -: col_length]};
assign pixels_row_14_22 = {data_out_rows[527*col_length-1 -: col_length]};
assign pixels_col_14_23 = {data_out_cols[528*col_length-1 -: col_length]};
assign pixels_row_14_23 = {data_out_rows[528*col_length-1 -: col_length]};
assign pixels_col_14_24 = {data_out_cols[529*col_length-1 -: col_length]};
assign pixels_row_14_24 = {data_out_rows[529*col_length-1 -: col_length]};
assign pixels_col_14_25 = {data_out_cols[530*col_length-1 -: col_length]};
assign pixels_row_14_25 = {data_out_rows[530*col_length-1 -: col_length]};
assign pixels_col_14_26 = {data_out_cols[531*col_length-1 -: col_length]};
assign pixels_row_14_26 = {data_out_rows[531*col_length-1 -: col_length]};
assign pixels_col_14_27 = {data_out_cols[532*col_length-1 -: col_length]};
assign pixels_row_14_27 = {data_out_rows[532*col_length-1 -: col_length]};
assign pixels_col_14_28 = {data_out_cols[533*col_length-1 -: col_length]};
assign pixels_row_14_28 = {data_out_rows[533*col_length-1 -: col_length]};
assign pixels_col_14_29 = {data_out_cols[534*col_length-1 -: col_length]};
assign pixels_row_14_29 = {data_out_rows[534*col_length-1 -: col_length]};
assign pixels_col_14_30 = {data_out_cols[535*col_length-1 -: col_length]};
assign pixels_row_14_30 = {data_out_rows[535*col_length-1 -: col_length]};
assign pixels_col_14_31 = {data_out_cols[536*col_length-1 -: col_length]};
assign pixels_row_14_31 = {data_out_rows[536*col_length-1 -: col_length]};
assign pixels_col_14_32 = {data_out_cols[537*col_length-1 -: col_length]};
assign pixels_row_14_32 = {data_out_rows[537*col_length-1 -: col_length]};
assign pixels_col_14_33 = {data_out_cols[538*col_length-1 -: col_length]};
assign pixels_row_14_33 = {data_out_rows[538*col_length-1 -: col_length]};
assign pixels_col_14_34 = {data_out_cols[539*col_length-1 -: col_length]};
assign pixels_row_14_34 = {data_out_rows[539*col_length-1 -: col_length]};
assign pixels_col_14_35 = {data_out_cols[540*col_length-1 -: col_length]};
assign pixels_row_14_35 = {data_out_rows[540*col_length-1 -: col_length]};
assign pixels_col_15_0 = {data_out_cols[541*col_length-1 -: col_length]};
assign pixels_row_15_0 = {data_out_rows[541*col_length-1 -: col_length]};
assign pixels_col_15_1 = {data_out_cols[542*col_length-1 -: col_length]};
assign pixels_row_15_1 = {data_out_rows[542*col_length-1 -: col_length]};
assign pixels_col_15_2 = {data_out_cols[543*col_length-1 -: col_length]};
assign pixels_row_15_2 = {data_out_rows[543*col_length-1 -: col_length]};
assign pixels_col_15_3 = {data_out_cols[544*col_length-1 -: col_length]};
assign pixels_row_15_3 = {data_out_rows[544*col_length-1 -: col_length]};
assign pixels_col_15_4 = {data_out_cols[545*col_length-1 -: col_length]};
assign pixels_row_15_4 = {data_out_rows[545*col_length-1 -: col_length]};
assign pixels_col_15_5 = {data_out_cols[546*col_length-1 -: col_length]};
assign pixels_row_15_5 = {data_out_rows[546*col_length-1 -: col_length]};
assign pixels_col_15_6 = {data_out_cols[547*col_length-1 -: col_length]};
assign pixels_row_15_6 = {data_out_rows[547*col_length-1 -: col_length]};
assign pixels_col_15_7 = {data_out_cols[548*col_length-1 -: col_length]};
assign pixels_row_15_7 = {data_out_rows[548*col_length-1 -: col_length]};
assign pixels_col_15_8 = {data_out_cols[549*col_length-1 -: col_length]};
assign pixels_row_15_8 = {data_out_rows[549*col_length-1 -: col_length]};
assign pixels_col_15_9 = {data_out_cols[550*col_length-1 -: col_length]};
assign pixels_row_15_9 = {data_out_rows[550*col_length-1 -: col_length]};
assign pixels_col_15_10 = {data_out_cols[551*col_length-1 -: col_length]};
assign pixels_row_15_10 = {data_out_rows[551*col_length-1 -: col_length]};
assign pixels_col_15_11 = {data_out_cols[552*col_length-1 -: col_length]};
assign pixels_row_15_11 = {data_out_rows[552*col_length-1 -: col_length]};
assign pixels_col_15_12 = {data_out_cols[553*col_length-1 -: col_length]};
assign pixels_row_15_12 = {data_out_rows[553*col_length-1 -: col_length]};
assign pixels_col_15_13 = {data_out_cols[554*col_length-1 -: col_length]};
assign pixels_row_15_13 = {data_out_rows[554*col_length-1 -: col_length]};
assign pixels_col_15_14 = {data_out_cols[555*col_length-1 -: col_length]};
assign pixels_row_15_14 = {data_out_rows[555*col_length-1 -: col_length]};
assign pixels_col_15_15 = {data_out_cols[556*col_length-1 -: col_length]};
assign pixels_row_15_15 = {data_out_rows[556*col_length-1 -: col_length]};
assign pixels_col_15_16 = {data_out_cols[557*col_length-1 -: col_length]};
assign pixels_row_15_16 = {data_out_rows[557*col_length-1 -: col_length]};
assign pixels_col_15_17 = {data_out_cols[558*col_length-1 -: col_length]};
assign pixels_row_15_17 = {data_out_rows[558*col_length-1 -: col_length]};
assign pixels_col_15_18 = {data_out_cols[559*col_length-1 -: col_length]};
assign pixels_row_15_18 = {data_out_rows[559*col_length-1 -: col_length]};
assign pixels_col_15_19 = {data_out_cols[560*col_length-1 -: col_length]};
assign pixels_row_15_19 = {data_out_rows[560*col_length-1 -: col_length]};
assign pixels_col_15_20 = {data_out_cols[561*col_length-1 -: col_length]};
assign pixels_row_15_20 = {data_out_rows[561*col_length-1 -: col_length]};
assign pixels_col_15_21 = {data_out_cols[562*col_length-1 -: col_length]};
assign pixels_row_15_21 = {data_out_rows[562*col_length-1 -: col_length]};
assign pixels_col_15_22 = {data_out_cols[563*col_length-1 -: col_length]};
assign pixels_row_15_22 = {data_out_rows[563*col_length-1 -: col_length]};
assign pixels_col_15_23 = {data_out_cols[564*col_length-1 -: col_length]};
assign pixels_row_15_23 = {data_out_rows[564*col_length-1 -: col_length]};
assign pixels_col_15_24 = {data_out_cols[565*col_length-1 -: col_length]};
assign pixels_row_15_24 = {data_out_rows[565*col_length-1 -: col_length]};
assign pixels_col_15_25 = {data_out_cols[566*col_length-1 -: col_length]};
assign pixels_row_15_25 = {data_out_rows[566*col_length-1 -: col_length]};
assign pixels_col_15_26 = {data_out_cols[567*col_length-1 -: col_length]};
assign pixels_row_15_26 = {data_out_rows[567*col_length-1 -: col_length]};
assign pixels_col_15_27 = {data_out_cols[568*col_length-1 -: col_length]};
assign pixels_row_15_27 = {data_out_rows[568*col_length-1 -: col_length]};
assign pixels_col_15_28 = {data_out_cols[569*col_length-1 -: col_length]};
assign pixels_row_15_28 = {data_out_rows[569*col_length-1 -: col_length]};
assign pixels_col_15_29 = {data_out_cols[570*col_length-1 -: col_length]};
assign pixels_row_15_29 = {data_out_rows[570*col_length-1 -: col_length]};
assign pixels_col_15_30 = {data_out_cols[571*col_length-1 -: col_length]};
assign pixels_row_15_30 = {data_out_rows[571*col_length-1 -: col_length]};
assign pixels_col_15_31 = {data_out_cols[572*col_length-1 -: col_length]};
assign pixels_row_15_31 = {data_out_rows[572*col_length-1 -: col_length]};
assign pixels_col_15_32 = {data_out_cols[573*col_length-1 -: col_length]};
assign pixels_row_15_32 = {data_out_rows[573*col_length-1 -: col_length]};
assign pixels_col_15_33 = {data_out_cols[574*col_length-1 -: col_length]};
assign pixels_row_15_33 = {data_out_rows[574*col_length-1 -: col_length]};
assign pixels_col_15_34 = {data_out_cols[575*col_length-1 -: col_length]};
assign pixels_row_15_34 = {data_out_rows[575*col_length-1 -: col_length]};
assign pixels_col_15_35 = {data_out_cols[576*col_length-1 -: col_length]};
assign pixels_row_15_35 = {data_out_rows[576*col_length-1 -: col_length]};
assign pixels_col_16_0 = {data_out_cols[577*col_length-1 -: col_length]};
assign pixels_row_16_0 = {data_out_rows[577*col_length-1 -: col_length]};
assign pixels_col_16_1 = {data_out_cols[578*col_length-1 -: col_length]};
assign pixels_row_16_1 = {data_out_rows[578*col_length-1 -: col_length]};
assign pixels_col_16_2 = {data_out_cols[579*col_length-1 -: col_length]};
assign pixels_row_16_2 = {data_out_rows[579*col_length-1 -: col_length]};
assign pixels_col_16_3 = {data_out_cols[580*col_length-1 -: col_length]};
assign pixels_row_16_3 = {data_out_rows[580*col_length-1 -: col_length]};
assign pixels_col_16_4 = {data_out_cols[581*col_length-1 -: col_length]};
assign pixels_row_16_4 = {data_out_rows[581*col_length-1 -: col_length]};
assign pixels_col_16_5 = {data_out_cols[582*col_length-1 -: col_length]};
assign pixels_row_16_5 = {data_out_rows[582*col_length-1 -: col_length]};
assign pixels_col_16_6 = {data_out_cols[583*col_length-1 -: col_length]};
assign pixels_row_16_6 = {data_out_rows[583*col_length-1 -: col_length]};
assign pixels_col_16_7 = {data_out_cols[584*col_length-1 -: col_length]};
assign pixels_row_16_7 = {data_out_rows[584*col_length-1 -: col_length]};
assign pixels_col_16_8 = {data_out_cols[585*col_length-1 -: col_length]};
assign pixels_row_16_8 = {data_out_rows[585*col_length-1 -: col_length]};
assign pixels_col_16_9 = {data_out_cols[586*col_length-1 -: col_length]};
assign pixels_row_16_9 = {data_out_rows[586*col_length-1 -: col_length]};
assign pixels_col_16_10 = {data_out_cols[587*col_length-1 -: col_length]};
assign pixels_row_16_10 = {data_out_rows[587*col_length-1 -: col_length]};
assign pixels_col_16_11 = {data_out_cols[588*col_length-1 -: col_length]};
assign pixels_row_16_11 = {data_out_rows[588*col_length-1 -: col_length]};
assign pixels_col_16_12 = {data_out_cols[589*col_length-1 -: col_length]};
assign pixels_row_16_12 = {data_out_rows[589*col_length-1 -: col_length]};
assign pixels_col_16_13 = {data_out_cols[590*col_length-1 -: col_length]};
assign pixels_row_16_13 = {data_out_rows[590*col_length-1 -: col_length]};
assign pixels_col_16_14 = {data_out_cols[591*col_length-1 -: col_length]};
assign pixels_row_16_14 = {data_out_rows[591*col_length-1 -: col_length]};
assign pixels_col_16_15 = {data_out_cols[592*col_length-1 -: col_length]};
assign pixels_row_16_15 = {data_out_rows[592*col_length-1 -: col_length]};
assign pixels_col_16_16 = {data_out_cols[593*col_length-1 -: col_length]};
assign pixels_row_16_16 = {data_out_rows[593*col_length-1 -: col_length]};
assign pixels_col_16_17 = {data_out_cols[594*col_length-1 -: col_length]};
assign pixels_row_16_17 = {data_out_rows[594*col_length-1 -: col_length]};
assign pixels_col_16_18 = {data_out_cols[595*col_length-1 -: col_length]};
assign pixels_row_16_18 = {data_out_rows[595*col_length-1 -: col_length]};
assign pixels_col_16_19 = {data_out_cols[596*col_length-1 -: col_length]};
assign pixels_row_16_19 = {data_out_rows[596*col_length-1 -: col_length]};
assign pixels_col_16_20 = {data_out_cols[597*col_length-1 -: col_length]};
assign pixels_row_16_20 = {data_out_rows[597*col_length-1 -: col_length]};
assign pixels_col_16_21 = {data_out_cols[598*col_length-1 -: col_length]};
assign pixels_row_16_21 = {data_out_rows[598*col_length-1 -: col_length]};
assign pixels_col_16_22 = {data_out_cols[599*col_length-1 -: col_length]};
assign pixels_row_16_22 = {data_out_rows[599*col_length-1 -: col_length]};
assign pixels_col_16_23 = {data_out_cols[600*col_length-1 -: col_length]};
assign pixels_row_16_23 = {data_out_rows[600*col_length-1 -: col_length]};
assign pixels_col_16_24 = {data_out_cols[601*col_length-1 -: col_length]};
assign pixels_row_16_24 = {data_out_rows[601*col_length-1 -: col_length]};
assign pixels_col_16_25 = {data_out_cols[602*col_length-1 -: col_length]};
assign pixels_row_16_25 = {data_out_rows[602*col_length-1 -: col_length]};
assign pixels_col_16_26 = {data_out_cols[603*col_length-1 -: col_length]};
assign pixels_row_16_26 = {data_out_rows[603*col_length-1 -: col_length]};
assign pixels_col_16_27 = {data_out_cols[604*col_length-1 -: col_length]};
assign pixels_row_16_27 = {data_out_rows[604*col_length-1 -: col_length]};
assign pixels_col_16_28 = {data_out_cols[605*col_length-1 -: col_length]};
assign pixels_row_16_28 = {data_out_rows[605*col_length-1 -: col_length]};
assign pixels_col_16_29 = {data_out_cols[606*col_length-1 -: col_length]};
assign pixels_row_16_29 = {data_out_rows[606*col_length-1 -: col_length]};
assign pixels_col_16_30 = {data_out_cols[607*col_length-1 -: col_length]};
assign pixels_row_16_30 = {data_out_rows[607*col_length-1 -: col_length]};
assign pixels_col_16_31 = {data_out_cols[608*col_length-1 -: col_length]};
assign pixels_row_16_31 = {data_out_rows[608*col_length-1 -: col_length]};
assign pixels_col_16_32 = {data_out_cols[609*col_length-1 -: col_length]};
assign pixels_row_16_32 = {data_out_rows[609*col_length-1 -: col_length]};
assign pixels_col_16_33 = {data_out_cols[610*col_length-1 -: col_length]};
assign pixels_row_16_33 = {data_out_rows[610*col_length-1 -: col_length]};
assign pixels_col_16_34 = {data_out_cols[611*col_length-1 -: col_length]};
assign pixels_row_16_34 = {data_out_rows[611*col_length-1 -: col_length]};
assign pixels_col_16_35 = {data_out_cols[612*col_length-1 -: col_length]};
assign pixels_row_16_35 = {data_out_rows[612*col_length-1 -: col_length]};
assign pixels_col_17_0 = {data_out_cols[613*col_length-1 -: col_length]};
assign pixels_row_17_0 = {data_out_rows[613*col_length-1 -: col_length]};
assign pixels_col_17_1 = {data_out_cols[614*col_length-1 -: col_length]};
assign pixels_row_17_1 = {data_out_rows[614*col_length-1 -: col_length]};
assign pixels_col_17_2 = {data_out_cols[615*col_length-1 -: col_length]};
assign pixels_row_17_2 = {data_out_rows[615*col_length-1 -: col_length]};
assign pixels_col_17_3 = {data_out_cols[616*col_length-1 -: col_length]};
assign pixels_row_17_3 = {data_out_rows[616*col_length-1 -: col_length]};
assign pixels_col_17_4 = {data_out_cols[617*col_length-1 -: col_length]};
assign pixels_row_17_4 = {data_out_rows[617*col_length-1 -: col_length]};
assign pixels_col_17_5 = {data_out_cols[618*col_length-1 -: col_length]};
assign pixels_row_17_5 = {data_out_rows[618*col_length-1 -: col_length]};
assign pixels_col_17_6 = {data_out_cols[619*col_length-1 -: col_length]};
assign pixels_row_17_6 = {data_out_rows[619*col_length-1 -: col_length]};
assign pixels_col_17_7 = {data_out_cols[620*col_length-1 -: col_length]};
assign pixels_row_17_7 = {data_out_rows[620*col_length-1 -: col_length]};
assign pixels_col_17_8 = {data_out_cols[621*col_length-1 -: col_length]};
assign pixels_row_17_8 = {data_out_rows[621*col_length-1 -: col_length]};
assign pixels_col_17_9 = {data_out_cols[622*col_length-1 -: col_length]};
assign pixels_row_17_9 = {data_out_rows[622*col_length-1 -: col_length]};
assign pixels_col_17_10 = {data_out_cols[623*col_length-1 -: col_length]};
assign pixels_row_17_10 = {data_out_rows[623*col_length-1 -: col_length]};
assign pixels_col_17_11 = {data_out_cols[624*col_length-1 -: col_length]};
assign pixels_row_17_11 = {data_out_rows[624*col_length-1 -: col_length]};
assign pixels_col_17_12 = {data_out_cols[625*col_length-1 -: col_length]};
assign pixels_row_17_12 = {data_out_rows[625*col_length-1 -: col_length]};
assign pixels_col_17_13 = {data_out_cols[626*col_length-1 -: col_length]};
assign pixels_row_17_13 = {data_out_rows[626*col_length-1 -: col_length]};
assign pixels_col_17_14 = {data_out_cols[627*col_length-1 -: col_length]};
assign pixels_row_17_14 = {data_out_rows[627*col_length-1 -: col_length]};
assign pixels_col_17_15 = {data_out_cols[628*col_length-1 -: col_length]};
assign pixels_row_17_15 = {data_out_rows[628*col_length-1 -: col_length]};
assign pixels_col_17_16 = {data_out_cols[629*col_length-1 -: col_length]};
assign pixels_row_17_16 = {data_out_rows[629*col_length-1 -: col_length]};
assign pixels_col_17_17 = {data_out_cols[630*col_length-1 -: col_length]};
assign pixels_row_17_17 = {data_out_rows[630*col_length-1 -: col_length]};
assign pixels_col_17_18 = {data_out_cols[631*col_length-1 -: col_length]};
assign pixels_row_17_18 = {data_out_rows[631*col_length-1 -: col_length]};
assign pixels_col_17_19 = {data_out_cols[632*col_length-1 -: col_length]};
assign pixels_row_17_19 = {data_out_rows[632*col_length-1 -: col_length]};
assign pixels_col_17_20 = {data_out_cols[633*col_length-1 -: col_length]};
assign pixels_row_17_20 = {data_out_rows[633*col_length-1 -: col_length]};
assign pixels_col_17_21 = {data_out_cols[634*col_length-1 -: col_length]};
assign pixels_row_17_21 = {data_out_rows[634*col_length-1 -: col_length]};
assign pixels_col_17_22 = {data_out_cols[635*col_length-1 -: col_length]};
assign pixels_row_17_22 = {data_out_rows[635*col_length-1 -: col_length]};
assign pixels_col_17_23 = {data_out_cols[636*col_length-1 -: col_length]};
assign pixels_row_17_23 = {data_out_rows[636*col_length-1 -: col_length]};
assign pixels_col_17_24 = {data_out_cols[637*col_length-1 -: col_length]};
assign pixels_row_17_24 = {data_out_rows[637*col_length-1 -: col_length]};
assign pixels_col_17_25 = {data_out_cols[638*col_length-1 -: col_length]};
assign pixels_row_17_25 = {data_out_rows[638*col_length-1 -: col_length]};
assign pixels_col_17_26 = {data_out_cols[639*col_length-1 -: col_length]};
assign pixels_row_17_26 = {data_out_rows[639*col_length-1 -: col_length]};
assign pixels_col_17_27 = {data_out_cols[640*col_length-1 -: col_length]};
assign pixels_row_17_27 = {data_out_rows[640*col_length-1 -: col_length]};
assign pixels_col_17_28 = {data_out_cols[641*col_length-1 -: col_length]};
assign pixels_row_17_28 = {data_out_rows[641*col_length-1 -: col_length]};
assign pixels_col_17_29 = {data_out_cols[642*col_length-1 -: col_length]};
assign pixels_row_17_29 = {data_out_rows[642*col_length-1 -: col_length]};
assign pixels_col_17_30 = {data_out_cols[643*col_length-1 -: col_length]};
assign pixels_row_17_30 = {data_out_rows[643*col_length-1 -: col_length]};
assign pixels_col_17_31 = {data_out_cols[644*col_length-1 -: col_length]};
assign pixels_row_17_31 = {data_out_rows[644*col_length-1 -: col_length]};
assign pixels_col_17_32 = {data_out_cols[645*col_length-1 -: col_length]};
assign pixels_row_17_32 = {data_out_rows[645*col_length-1 -: col_length]};
assign pixels_col_17_33 = {data_out_cols[646*col_length-1 -: col_length]};
assign pixels_row_17_33 = {data_out_rows[646*col_length-1 -: col_length]};
assign pixels_col_17_34 = {data_out_cols[647*col_length-1 -: col_length]};
assign pixels_row_17_34 = {data_out_rows[647*col_length-1 -: col_length]};
assign pixels_col_17_35 = {data_out_cols[648*col_length-1 -: col_length]};
assign pixels_row_17_35 = {data_out_rows[648*col_length-1 -: col_length]};
assign pixels_col_18_0 = {data_out_cols[649*col_length-1 -: col_length]};
assign pixels_row_18_0 = {data_out_rows[649*col_length-1 -: col_length]};
assign pixels_col_18_1 = {data_out_cols[650*col_length-1 -: col_length]};
assign pixels_row_18_1 = {data_out_rows[650*col_length-1 -: col_length]};
assign pixels_col_18_2 = {data_out_cols[651*col_length-1 -: col_length]};
assign pixels_row_18_2 = {data_out_rows[651*col_length-1 -: col_length]};
assign pixels_col_18_3 = {data_out_cols[652*col_length-1 -: col_length]};
assign pixels_row_18_3 = {data_out_rows[652*col_length-1 -: col_length]};
assign pixels_col_18_4 = {data_out_cols[653*col_length-1 -: col_length]};
assign pixels_row_18_4 = {data_out_rows[653*col_length-1 -: col_length]};
assign pixels_col_18_5 = {data_out_cols[654*col_length-1 -: col_length]};
assign pixels_row_18_5 = {data_out_rows[654*col_length-1 -: col_length]};
assign pixels_col_18_6 = {data_out_cols[655*col_length-1 -: col_length]};
assign pixels_row_18_6 = {data_out_rows[655*col_length-1 -: col_length]};
assign pixels_col_18_7 = {data_out_cols[656*col_length-1 -: col_length]};
assign pixels_row_18_7 = {data_out_rows[656*col_length-1 -: col_length]};
assign pixels_col_18_8 = {data_out_cols[657*col_length-1 -: col_length]};
assign pixels_row_18_8 = {data_out_rows[657*col_length-1 -: col_length]};
assign pixels_col_18_9 = {data_out_cols[658*col_length-1 -: col_length]};
assign pixels_row_18_9 = {data_out_rows[658*col_length-1 -: col_length]};
assign pixels_col_18_10 = {data_out_cols[659*col_length-1 -: col_length]};
assign pixels_row_18_10 = {data_out_rows[659*col_length-1 -: col_length]};
assign pixels_col_18_11 = {data_out_cols[660*col_length-1 -: col_length]};
assign pixels_row_18_11 = {data_out_rows[660*col_length-1 -: col_length]};
assign pixels_col_18_12 = {data_out_cols[661*col_length-1 -: col_length]};
assign pixels_row_18_12 = {data_out_rows[661*col_length-1 -: col_length]};
assign pixels_col_18_13 = {data_out_cols[662*col_length-1 -: col_length]};
assign pixels_row_18_13 = {data_out_rows[662*col_length-1 -: col_length]};
assign pixels_col_18_14 = {data_out_cols[663*col_length-1 -: col_length]};
assign pixels_row_18_14 = {data_out_rows[663*col_length-1 -: col_length]};
assign pixels_col_18_15 = {data_out_cols[664*col_length-1 -: col_length]};
assign pixels_row_18_15 = {data_out_rows[664*col_length-1 -: col_length]};
assign pixels_col_18_16 = {data_out_cols[665*col_length-1 -: col_length]};
assign pixels_row_18_16 = {data_out_rows[665*col_length-1 -: col_length]};
assign pixels_col_18_17 = {data_out_cols[666*col_length-1 -: col_length]};
assign pixels_row_18_17 = {data_out_rows[666*col_length-1 -: col_length]};
assign pixels_col_18_18 = {data_out_cols[667*col_length-1 -: col_length]};
assign pixels_row_18_18 = {data_out_rows[667*col_length-1 -: col_length]};
assign pixels_col_18_19 = {data_out_cols[668*col_length-1 -: col_length]};
assign pixels_row_18_19 = {data_out_rows[668*col_length-1 -: col_length]};
assign pixels_col_18_20 = {data_out_cols[669*col_length-1 -: col_length]};
assign pixels_row_18_20 = {data_out_rows[669*col_length-1 -: col_length]};
assign pixels_col_18_21 = {data_out_cols[670*col_length-1 -: col_length]};
assign pixels_row_18_21 = {data_out_rows[670*col_length-1 -: col_length]};
assign pixels_col_18_22 = {data_out_cols[671*col_length-1 -: col_length]};
assign pixels_row_18_22 = {data_out_rows[671*col_length-1 -: col_length]};
assign pixels_col_18_23 = {data_out_cols[672*col_length-1 -: col_length]};
assign pixels_row_18_23 = {data_out_rows[672*col_length-1 -: col_length]};
assign pixels_col_18_24 = {data_out_cols[673*col_length-1 -: col_length]};
assign pixels_row_18_24 = {data_out_rows[673*col_length-1 -: col_length]};
assign pixels_col_18_25 = {data_out_cols[674*col_length-1 -: col_length]};
assign pixels_row_18_25 = {data_out_rows[674*col_length-1 -: col_length]};
assign pixels_col_18_26 = {data_out_cols[675*col_length-1 -: col_length]};
assign pixels_row_18_26 = {data_out_rows[675*col_length-1 -: col_length]};
assign pixels_col_18_27 = {data_out_cols[676*col_length-1 -: col_length]};
assign pixels_row_18_27 = {data_out_rows[676*col_length-1 -: col_length]};
assign pixels_col_18_28 = {data_out_cols[677*col_length-1 -: col_length]};
assign pixels_row_18_28 = {data_out_rows[677*col_length-1 -: col_length]};
assign pixels_col_18_29 = {data_out_cols[678*col_length-1 -: col_length]};
assign pixels_row_18_29 = {data_out_rows[678*col_length-1 -: col_length]};
assign pixels_col_18_30 = {data_out_cols[679*col_length-1 -: col_length]};
assign pixels_row_18_30 = {data_out_rows[679*col_length-1 -: col_length]};
assign pixels_col_18_31 = {data_out_cols[680*col_length-1 -: col_length]};
assign pixels_row_18_31 = {data_out_rows[680*col_length-1 -: col_length]};
assign pixels_col_18_32 = {data_out_cols[681*col_length-1 -: col_length]};
assign pixels_row_18_32 = {data_out_rows[681*col_length-1 -: col_length]};
assign pixels_col_18_33 = {data_out_cols[682*col_length-1 -: col_length]};
assign pixels_row_18_33 = {data_out_rows[682*col_length-1 -: col_length]};
assign pixels_col_18_34 = {data_out_cols[683*col_length-1 -: col_length]};
assign pixels_row_18_34 = {data_out_rows[683*col_length-1 -: col_length]};
assign pixels_col_18_35 = {data_out_cols[684*col_length-1 -: col_length]};
assign pixels_row_18_35 = {data_out_rows[684*col_length-1 -: col_length]};
assign pixels_col_19_0 = {data_out_cols[685*col_length-1 -: col_length]};
assign pixels_row_19_0 = {data_out_rows[685*col_length-1 -: col_length]};
assign pixels_col_19_1 = {data_out_cols[686*col_length-1 -: col_length]};
assign pixels_row_19_1 = {data_out_rows[686*col_length-1 -: col_length]};
assign pixels_col_19_2 = {data_out_cols[687*col_length-1 -: col_length]};
assign pixels_row_19_2 = {data_out_rows[687*col_length-1 -: col_length]};
assign pixels_col_19_3 = {data_out_cols[688*col_length-1 -: col_length]};
assign pixels_row_19_3 = {data_out_rows[688*col_length-1 -: col_length]};
assign pixels_col_19_4 = {data_out_cols[689*col_length-1 -: col_length]};
assign pixels_row_19_4 = {data_out_rows[689*col_length-1 -: col_length]};
assign pixels_col_19_5 = {data_out_cols[690*col_length-1 -: col_length]};
assign pixels_row_19_5 = {data_out_rows[690*col_length-1 -: col_length]};
assign pixels_col_19_6 = {data_out_cols[691*col_length-1 -: col_length]};
assign pixels_row_19_6 = {data_out_rows[691*col_length-1 -: col_length]};
assign pixels_col_19_7 = {data_out_cols[692*col_length-1 -: col_length]};
assign pixels_row_19_7 = {data_out_rows[692*col_length-1 -: col_length]};
assign pixels_col_19_8 = {data_out_cols[693*col_length-1 -: col_length]};
assign pixels_row_19_8 = {data_out_rows[693*col_length-1 -: col_length]};
assign pixels_col_19_9 = {data_out_cols[694*col_length-1 -: col_length]};
assign pixels_row_19_9 = {data_out_rows[694*col_length-1 -: col_length]};
assign pixels_col_19_10 = {data_out_cols[695*col_length-1 -: col_length]};
assign pixels_row_19_10 = {data_out_rows[695*col_length-1 -: col_length]};
assign pixels_col_19_11 = {data_out_cols[696*col_length-1 -: col_length]};
assign pixels_row_19_11 = {data_out_rows[696*col_length-1 -: col_length]};
assign pixels_col_19_12 = {data_out_cols[697*col_length-1 -: col_length]};
assign pixels_row_19_12 = {data_out_rows[697*col_length-1 -: col_length]};
assign pixels_col_19_13 = {data_out_cols[698*col_length-1 -: col_length]};
assign pixels_row_19_13 = {data_out_rows[698*col_length-1 -: col_length]};
assign pixels_col_19_14 = {data_out_cols[699*col_length-1 -: col_length]};
assign pixels_row_19_14 = {data_out_rows[699*col_length-1 -: col_length]};
assign pixels_col_19_15 = {data_out_cols[700*col_length-1 -: col_length]};
assign pixels_row_19_15 = {data_out_rows[700*col_length-1 -: col_length]};
assign pixels_col_19_16 = {data_out_cols[701*col_length-1 -: col_length]};
assign pixels_row_19_16 = {data_out_rows[701*col_length-1 -: col_length]};
assign pixels_col_19_17 = {data_out_cols[702*col_length-1 -: col_length]};
assign pixels_row_19_17 = {data_out_rows[702*col_length-1 -: col_length]};
assign pixels_col_19_18 = {data_out_cols[703*col_length-1 -: col_length]};
assign pixels_row_19_18 = {data_out_rows[703*col_length-1 -: col_length]};
assign pixels_col_19_19 = {data_out_cols[704*col_length-1 -: col_length]};
assign pixels_row_19_19 = {data_out_rows[704*col_length-1 -: col_length]};
assign pixels_col_19_20 = {data_out_cols[705*col_length-1 -: col_length]};
assign pixels_row_19_20 = {data_out_rows[705*col_length-1 -: col_length]};
assign pixels_col_19_21 = {data_out_cols[706*col_length-1 -: col_length]};
assign pixels_row_19_21 = {data_out_rows[706*col_length-1 -: col_length]};
assign pixels_col_19_22 = {data_out_cols[707*col_length-1 -: col_length]};
assign pixels_row_19_22 = {data_out_rows[707*col_length-1 -: col_length]};
assign pixels_col_19_23 = {data_out_cols[708*col_length-1 -: col_length]};
assign pixels_row_19_23 = {data_out_rows[708*col_length-1 -: col_length]};
assign pixels_col_19_24 = {data_out_cols[709*col_length-1 -: col_length]};
assign pixels_row_19_24 = {data_out_rows[709*col_length-1 -: col_length]};
assign pixels_col_19_25 = {data_out_cols[710*col_length-1 -: col_length]};
assign pixels_row_19_25 = {data_out_rows[710*col_length-1 -: col_length]};
assign pixels_col_19_26 = {data_out_cols[711*col_length-1 -: col_length]};
assign pixels_row_19_26 = {data_out_rows[711*col_length-1 -: col_length]};
assign pixels_col_19_27 = {data_out_cols[712*col_length-1 -: col_length]};
assign pixels_row_19_27 = {data_out_rows[712*col_length-1 -: col_length]};
assign pixels_col_19_28 = {data_out_cols[713*col_length-1 -: col_length]};
assign pixels_row_19_28 = {data_out_rows[713*col_length-1 -: col_length]};
assign pixels_col_19_29 = {data_out_cols[714*col_length-1 -: col_length]};
assign pixels_row_19_29 = {data_out_rows[714*col_length-1 -: col_length]};
assign pixels_col_19_30 = {data_out_cols[715*col_length-1 -: col_length]};
assign pixels_row_19_30 = {data_out_rows[715*col_length-1 -: col_length]};
assign pixels_col_19_31 = {data_out_cols[716*col_length-1 -: col_length]};
assign pixels_row_19_31 = {data_out_rows[716*col_length-1 -: col_length]};
assign pixels_col_19_32 = {data_out_cols[717*col_length-1 -: col_length]};
assign pixels_row_19_32 = {data_out_rows[717*col_length-1 -: col_length]};
assign pixels_col_19_33 = {data_out_cols[718*col_length-1 -: col_length]};
assign pixels_row_19_33 = {data_out_rows[718*col_length-1 -: col_length]};
assign pixels_col_19_34 = {data_out_cols[719*col_length-1 -: col_length]};
assign pixels_row_19_34 = {data_out_rows[719*col_length-1 -: col_length]};
assign pixels_col_19_35 = {data_out_cols[720*col_length-1 -: col_length]};
assign pixels_row_19_35 = {data_out_rows[720*col_length-1 -: col_length]};
assign pixels_col_20_0 = {data_out_cols[721*col_length-1 -: col_length]};
assign pixels_row_20_0 = {data_out_rows[721*col_length-1 -: col_length]};
assign pixels_col_20_1 = {data_out_cols[722*col_length-1 -: col_length]};
assign pixels_row_20_1 = {data_out_rows[722*col_length-1 -: col_length]};
assign pixels_col_20_2 = {data_out_cols[723*col_length-1 -: col_length]};
assign pixels_row_20_2 = {data_out_rows[723*col_length-1 -: col_length]};
assign pixels_col_20_3 = {data_out_cols[724*col_length-1 -: col_length]};
assign pixels_row_20_3 = {data_out_rows[724*col_length-1 -: col_length]};
assign pixels_col_20_4 = {data_out_cols[725*col_length-1 -: col_length]};
assign pixels_row_20_4 = {data_out_rows[725*col_length-1 -: col_length]};
assign pixels_col_20_5 = {data_out_cols[726*col_length-1 -: col_length]};
assign pixels_row_20_5 = {data_out_rows[726*col_length-1 -: col_length]};
assign pixels_col_20_6 = {data_out_cols[727*col_length-1 -: col_length]};
assign pixels_row_20_6 = {data_out_rows[727*col_length-1 -: col_length]};
assign pixels_col_20_7 = {data_out_cols[728*col_length-1 -: col_length]};
assign pixels_row_20_7 = {data_out_rows[728*col_length-1 -: col_length]};
assign pixels_col_20_8 = {data_out_cols[729*col_length-1 -: col_length]};
assign pixels_row_20_8 = {data_out_rows[729*col_length-1 -: col_length]};
assign pixels_col_20_9 = {data_out_cols[730*col_length-1 -: col_length]};
assign pixels_row_20_9 = {data_out_rows[730*col_length-1 -: col_length]};
assign pixels_col_20_10 = {data_out_cols[731*col_length-1 -: col_length]};
assign pixels_row_20_10 = {data_out_rows[731*col_length-1 -: col_length]};
assign pixels_col_20_11 = {data_out_cols[732*col_length-1 -: col_length]};
assign pixels_row_20_11 = {data_out_rows[732*col_length-1 -: col_length]};
assign pixels_col_20_12 = {data_out_cols[733*col_length-1 -: col_length]};
assign pixels_row_20_12 = {data_out_rows[733*col_length-1 -: col_length]};
assign pixels_col_20_13 = {data_out_cols[734*col_length-1 -: col_length]};
assign pixels_row_20_13 = {data_out_rows[734*col_length-1 -: col_length]};
assign pixels_col_20_14 = {data_out_cols[735*col_length-1 -: col_length]};
assign pixels_row_20_14 = {data_out_rows[735*col_length-1 -: col_length]};
assign pixels_col_20_15 = {data_out_cols[736*col_length-1 -: col_length]};
assign pixels_row_20_15 = {data_out_rows[736*col_length-1 -: col_length]};
assign pixels_col_20_16 = {data_out_cols[737*col_length-1 -: col_length]};
assign pixels_row_20_16 = {data_out_rows[737*col_length-1 -: col_length]};
assign pixels_col_20_17 = {data_out_cols[738*col_length-1 -: col_length]};
assign pixels_row_20_17 = {data_out_rows[738*col_length-1 -: col_length]};
assign pixels_col_20_18 = {data_out_cols[739*col_length-1 -: col_length]};
assign pixels_row_20_18 = {data_out_rows[739*col_length-1 -: col_length]};
assign pixels_col_20_19 = {data_out_cols[740*col_length-1 -: col_length]};
assign pixels_row_20_19 = {data_out_rows[740*col_length-1 -: col_length]};
assign pixels_col_20_20 = {data_out_cols[741*col_length-1 -: col_length]};
assign pixels_row_20_20 = {data_out_rows[741*col_length-1 -: col_length]};
assign pixels_col_20_21 = {data_out_cols[742*col_length-1 -: col_length]};
assign pixels_row_20_21 = {data_out_rows[742*col_length-1 -: col_length]};
assign pixels_col_20_22 = {data_out_cols[743*col_length-1 -: col_length]};
assign pixels_row_20_22 = {data_out_rows[743*col_length-1 -: col_length]};
assign pixels_col_20_23 = {data_out_cols[744*col_length-1 -: col_length]};
assign pixels_row_20_23 = {data_out_rows[744*col_length-1 -: col_length]};
assign pixels_col_20_24 = {data_out_cols[745*col_length-1 -: col_length]};
assign pixels_row_20_24 = {data_out_rows[745*col_length-1 -: col_length]};
assign pixels_col_20_25 = {data_out_cols[746*col_length-1 -: col_length]};
assign pixels_row_20_25 = {data_out_rows[746*col_length-1 -: col_length]};
assign pixels_col_20_26 = {data_out_cols[747*col_length-1 -: col_length]};
assign pixels_row_20_26 = {data_out_rows[747*col_length-1 -: col_length]};
assign pixels_col_20_27 = {data_out_cols[748*col_length-1 -: col_length]};
assign pixels_row_20_27 = {data_out_rows[748*col_length-1 -: col_length]};
assign pixels_col_20_28 = {data_out_cols[749*col_length-1 -: col_length]};
assign pixels_row_20_28 = {data_out_rows[749*col_length-1 -: col_length]};
assign pixels_col_20_29 = {data_out_cols[750*col_length-1 -: col_length]};
assign pixels_row_20_29 = {data_out_rows[750*col_length-1 -: col_length]};
assign pixels_col_20_30 = {data_out_cols[751*col_length-1 -: col_length]};
assign pixels_row_20_30 = {data_out_rows[751*col_length-1 -: col_length]};
assign pixels_col_20_31 = {data_out_cols[752*col_length-1 -: col_length]};
assign pixels_row_20_31 = {data_out_rows[752*col_length-1 -: col_length]};
assign pixels_col_20_32 = {data_out_cols[753*col_length-1 -: col_length]};
assign pixels_row_20_32 = {data_out_rows[753*col_length-1 -: col_length]};
assign pixels_col_20_33 = {data_out_cols[754*col_length-1 -: col_length]};
assign pixels_row_20_33 = {data_out_rows[754*col_length-1 -: col_length]};
assign pixels_col_20_34 = {data_out_cols[755*col_length-1 -: col_length]};
assign pixels_row_20_34 = {data_out_rows[755*col_length-1 -: col_length]};
assign pixels_col_20_35 = {data_out_cols[756*col_length-1 -: col_length]};
assign pixels_row_20_35 = {data_out_rows[756*col_length-1 -: col_length]};
assign pixels_col_21_0 = {data_out_cols[757*col_length-1 -: col_length]};
assign pixels_row_21_0 = {data_out_rows[757*col_length-1 -: col_length]};
assign pixels_col_21_1 = {data_out_cols[758*col_length-1 -: col_length]};
assign pixels_row_21_1 = {data_out_rows[758*col_length-1 -: col_length]};
assign pixels_col_21_2 = {data_out_cols[759*col_length-1 -: col_length]};
assign pixels_row_21_2 = {data_out_rows[759*col_length-1 -: col_length]};
assign pixels_col_21_3 = {data_out_cols[760*col_length-1 -: col_length]};
assign pixels_row_21_3 = {data_out_rows[760*col_length-1 -: col_length]};
assign pixels_col_21_4 = {data_out_cols[761*col_length-1 -: col_length]};
assign pixels_row_21_4 = {data_out_rows[761*col_length-1 -: col_length]};
assign pixels_col_21_5 = {data_out_cols[762*col_length-1 -: col_length]};
assign pixels_row_21_5 = {data_out_rows[762*col_length-1 -: col_length]};
assign pixels_col_21_6 = {data_out_cols[763*col_length-1 -: col_length]};
assign pixels_row_21_6 = {data_out_rows[763*col_length-1 -: col_length]};
assign pixels_col_21_7 = {data_out_cols[764*col_length-1 -: col_length]};
assign pixels_row_21_7 = {data_out_rows[764*col_length-1 -: col_length]};
assign pixels_col_21_8 = {data_out_cols[765*col_length-1 -: col_length]};
assign pixels_row_21_8 = {data_out_rows[765*col_length-1 -: col_length]};
assign pixels_col_21_9 = {data_out_cols[766*col_length-1 -: col_length]};
assign pixels_row_21_9 = {data_out_rows[766*col_length-1 -: col_length]};
assign pixels_col_21_10 = {data_out_cols[767*col_length-1 -: col_length]};
assign pixels_row_21_10 = {data_out_rows[767*col_length-1 -: col_length]};
assign pixels_col_21_11 = {data_out_cols[768*col_length-1 -: col_length]};
assign pixels_row_21_11 = {data_out_rows[768*col_length-1 -: col_length]};
assign pixels_col_21_12 = {data_out_cols[769*col_length-1 -: col_length]};
assign pixels_row_21_12 = {data_out_rows[769*col_length-1 -: col_length]};
assign pixels_col_21_13 = {data_out_cols[770*col_length-1 -: col_length]};
assign pixels_row_21_13 = {data_out_rows[770*col_length-1 -: col_length]};
assign pixels_col_21_14 = {data_out_cols[771*col_length-1 -: col_length]};
assign pixels_row_21_14 = {data_out_rows[771*col_length-1 -: col_length]};
assign pixels_col_21_15 = {data_out_cols[772*col_length-1 -: col_length]};
assign pixels_row_21_15 = {data_out_rows[772*col_length-1 -: col_length]};
assign pixels_col_21_16 = {data_out_cols[773*col_length-1 -: col_length]};
assign pixels_row_21_16 = {data_out_rows[773*col_length-1 -: col_length]};
assign pixels_col_21_17 = {data_out_cols[774*col_length-1 -: col_length]};
assign pixels_row_21_17 = {data_out_rows[774*col_length-1 -: col_length]};
assign pixels_col_21_18 = {data_out_cols[775*col_length-1 -: col_length]};
assign pixels_row_21_18 = {data_out_rows[775*col_length-1 -: col_length]};
assign pixels_col_21_19 = {data_out_cols[776*col_length-1 -: col_length]};
assign pixels_row_21_19 = {data_out_rows[776*col_length-1 -: col_length]};
assign pixels_col_21_20 = {data_out_cols[777*col_length-1 -: col_length]};
assign pixels_row_21_20 = {data_out_rows[777*col_length-1 -: col_length]};
assign pixels_col_21_21 = {data_out_cols[778*col_length-1 -: col_length]};
assign pixels_row_21_21 = {data_out_rows[778*col_length-1 -: col_length]};
assign pixels_col_21_22 = {data_out_cols[779*col_length-1 -: col_length]};
assign pixels_row_21_22 = {data_out_rows[779*col_length-1 -: col_length]};
assign pixels_col_21_23 = {data_out_cols[780*col_length-1 -: col_length]};
assign pixels_row_21_23 = {data_out_rows[780*col_length-1 -: col_length]};
assign pixels_col_21_24 = {data_out_cols[781*col_length-1 -: col_length]};
assign pixels_row_21_24 = {data_out_rows[781*col_length-1 -: col_length]};
assign pixels_col_21_25 = {data_out_cols[782*col_length-1 -: col_length]};
assign pixels_row_21_25 = {data_out_rows[782*col_length-1 -: col_length]};
assign pixels_col_21_26 = {data_out_cols[783*col_length-1 -: col_length]};
assign pixels_row_21_26 = {data_out_rows[783*col_length-1 -: col_length]};
assign pixels_col_21_27 = {data_out_cols[784*col_length-1 -: col_length]};
assign pixels_row_21_27 = {data_out_rows[784*col_length-1 -: col_length]};
assign pixels_col_21_28 = {data_out_cols[785*col_length-1 -: col_length]};
assign pixels_row_21_28 = {data_out_rows[785*col_length-1 -: col_length]};
assign pixels_col_21_29 = {data_out_cols[786*col_length-1 -: col_length]};
assign pixels_row_21_29 = {data_out_rows[786*col_length-1 -: col_length]};
assign pixels_col_21_30 = {data_out_cols[787*col_length-1 -: col_length]};
assign pixels_row_21_30 = {data_out_rows[787*col_length-1 -: col_length]};
assign pixels_col_21_31 = {data_out_cols[788*col_length-1 -: col_length]};
assign pixels_row_21_31 = {data_out_rows[788*col_length-1 -: col_length]};
assign pixels_col_21_32 = {data_out_cols[789*col_length-1 -: col_length]};
assign pixels_row_21_32 = {data_out_rows[789*col_length-1 -: col_length]};
assign pixels_col_21_33 = {data_out_cols[790*col_length-1 -: col_length]};
assign pixels_row_21_33 = {data_out_rows[790*col_length-1 -: col_length]};
assign pixels_col_21_34 = {data_out_cols[791*col_length-1 -: col_length]};
assign pixels_row_21_34 = {data_out_rows[791*col_length-1 -: col_length]};
assign pixels_col_21_35 = {data_out_cols[792*col_length-1 -: col_length]};
assign pixels_row_21_35 = {data_out_rows[792*col_length-1 -: col_length]};
assign pixels_col_22_0 = {data_out_cols[793*col_length-1 -: col_length]};
assign pixels_row_22_0 = {data_out_rows[793*col_length-1 -: col_length]};
assign pixels_col_22_1 = {data_out_cols[794*col_length-1 -: col_length]};
assign pixels_row_22_1 = {data_out_rows[794*col_length-1 -: col_length]};
assign pixels_col_22_2 = {data_out_cols[795*col_length-1 -: col_length]};
assign pixels_row_22_2 = {data_out_rows[795*col_length-1 -: col_length]};
assign pixels_col_22_3 = {data_out_cols[796*col_length-1 -: col_length]};
assign pixels_row_22_3 = {data_out_rows[796*col_length-1 -: col_length]};
assign pixels_col_22_4 = {data_out_cols[797*col_length-1 -: col_length]};
assign pixels_row_22_4 = {data_out_rows[797*col_length-1 -: col_length]};
assign pixels_col_22_5 = {data_out_cols[798*col_length-1 -: col_length]};
assign pixels_row_22_5 = {data_out_rows[798*col_length-1 -: col_length]};
assign pixels_col_22_6 = {data_out_cols[799*col_length-1 -: col_length]};
assign pixels_row_22_6 = {data_out_rows[799*col_length-1 -: col_length]};
assign pixels_col_22_7 = {data_out_cols[800*col_length-1 -: col_length]};
assign pixels_row_22_7 = {data_out_rows[800*col_length-1 -: col_length]};
assign pixels_col_22_8 = {data_out_cols[801*col_length-1 -: col_length]};
assign pixels_row_22_8 = {data_out_rows[801*col_length-1 -: col_length]};
assign pixels_col_22_9 = {data_out_cols[802*col_length-1 -: col_length]};
assign pixels_row_22_9 = {data_out_rows[802*col_length-1 -: col_length]};
assign pixels_col_22_10 = {data_out_cols[803*col_length-1 -: col_length]};
assign pixels_row_22_10 = {data_out_rows[803*col_length-1 -: col_length]};
assign pixels_col_22_11 = {data_out_cols[804*col_length-1 -: col_length]};
assign pixels_row_22_11 = {data_out_rows[804*col_length-1 -: col_length]};
assign pixels_col_22_12 = {data_out_cols[805*col_length-1 -: col_length]};
assign pixels_row_22_12 = {data_out_rows[805*col_length-1 -: col_length]};
assign pixels_col_22_13 = {data_out_cols[806*col_length-1 -: col_length]};
assign pixels_row_22_13 = {data_out_rows[806*col_length-1 -: col_length]};
assign pixels_col_22_14 = {data_out_cols[807*col_length-1 -: col_length]};
assign pixels_row_22_14 = {data_out_rows[807*col_length-1 -: col_length]};
assign pixels_col_22_15 = {data_out_cols[808*col_length-1 -: col_length]};
assign pixels_row_22_15 = {data_out_rows[808*col_length-1 -: col_length]};
assign pixels_col_22_16 = {data_out_cols[809*col_length-1 -: col_length]};
assign pixels_row_22_16 = {data_out_rows[809*col_length-1 -: col_length]};
assign pixels_col_22_17 = {data_out_cols[810*col_length-1 -: col_length]};
assign pixels_row_22_17 = {data_out_rows[810*col_length-1 -: col_length]};
assign pixels_col_22_18 = {data_out_cols[811*col_length-1 -: col_length]};
assign pixels_row_22_18 = {data_out_rows[811*col_length-1 -: col_length]};
assign pixels_col_22_19 = {data_out_cols[812*col_length-1 -: col_length]};
assign pixels_row_22_19 = {data_out_rows[812*col_length-1 -: col_length]};
assign pixels_col_22_20 = {data_out_cols[813*col_length-1 -: col_length]};
assign pixels_row_22_20 = {data_out_rows[813*col_length-1 -: col_length]};
assign pixels_col_22_21 = {data_out_cols[814*col_length-1 -: col_length]};
assign pixels_row_22_21 = {data_out_rows[814*col_length-1 -: col_length]};
assign pixels_col_22_22 = {data_out_cols[815*col_length-1 -: col_length]};
assign pixels_row_22_22 = {data_out_rows[815*col_length-1 -: col_length]};
assign pixels_col_22_23 = {data_out_cols[816*col_length-1 -: col_length]};
assign pixels_row_22_23 = {data_out_rows[816*col_length-1 -: col_length]};
assign pixels_col_22_24 = {data_out_cols[817*col_length-1 -: col_length]};
assign pixels_row_22_24 = {data_out_rows[817*col_length-1 -: col_length]};
assign pixels_col_22_25 = {data_out_cols[818*col_length-1 -: col_length]};
assign pixels_row_22_25 = {data_out_rows[818*col_length-1 -: col_length]};
assign pixels_col_22_26 = {data_out_cols[819*col_length-1 -: col_length]};
assign pixels_row_22_26 = {data_out_rows[819*col_length-1 -: col_length]};
assign pixels_col_22_27 = {data_out_cols[820*col_length-1 -: col_length]};
assign pixels_row_22_27 = {data_out_rows[820*col_length-1 -: col_length]};
assign pixels_col_22_28 = {data_out_cols[821*col_length-1 -: col_length]};
assign pixels_row_22_28 = {data_out_rows[821*col_length-1 -: col_length]};
assign pixels_col_22_29 = {data_out_cols[822*col_length-1 -: col_length]};
assign pixels_row_22_29 = {data_out_rows[822*col_length-1 -: col_length]};
assign pixels_col_22_30 = {data_out_cols[823*col_length-1 -: col_length]};
assign pixels_row_22_30 = {data_out_rows[823*col_length-1 -: col_length]};
assign pixels_col_22_31 = {data_out_cols[824*col_length-1 -: col_length]};
assign pixels_row_22_31 = {data_out_rows[824*col_length-1 -: col_length]};
assign pixels_col_22_32 = {data_out_cols[825*col_length-1 -: col_length]};
assign pixels_row_22_32 = {data_out_rows[825*col_length-1 -: col_length]};
assign pixels_col_22_33 = {data_out_cols[826*col_length-1 -: col_length]};
assign pixels_row_22_33 = {data_out_rows[826*col_length-1 -: col_length]};
assign pixels_col_22_34 = {data_out_cols[827*col_length-1 -: col_length]};
assign pixels_row_22_34 = {data_out_rows[827*col_length-1 -: col_length]};
assign pixels_col_22_35 = {data_out_cols[828*col_length-1 -: col_length]};
assign pixels_row_22_35 = {data_out_rows[828*col_length-1 -: col_length]};
assign pixels_col_23_0 = {data_out_cols[829*col_length-1 -: col_length]};
assign pixels_row_23_0 = {data_out_rows[829*col_length-1 -: col_length]};
assign pixels_col_23_1 = {data_out_cols[830*col_length-1 -: col_length]};
assign pixels_row_23_1 = {data_out_rows[830*col_length-1 -: col_length]};
assign pixels_col_23_2 = {data_out_cols[831*col_length-1 -: col_length]};
assign pixels_row_23_2 = {data_out_rows[831*col_length-1 -: col_length]};
assign pixels_col_23_3 = {data_out_cols[832*col_length-1 -: col_length]};
assign pixels_row_23_3 = {data_out_rows[832*col_length-1 -: col_length]};
assign pixels_col_23_4 = {data_out_cols[833*col_length-1 -: col_length]};
assign pixels_row_23_4 = {data_out_rows[833*col_length-1 -: col_length]};
assign pixels_col_23_5 = {data_out_cols[834*col_length-1 -: col_length]};
assign pixels_row_23_5 = {data_out_rows[834*col_length-1 -: col_length]};
assign pixels_col_23_6 = {data_out_cols[835*col_length-1 -: col_length]};
assign pixels_row_23_6 = {data_out_rows[835*col_length-1 -: col_length]};
assign pixels_col_23_7 = {data_out_cols[836*col_length-1 -: col_length]};
assign pixels_row_23_7 = {data_out_rows[836*col_length-1 -: col_length]};
assign pixels_col_23_8 = {data_out_cols[837*col_length-1 -: col_length]};
assign pixels_row_23_8 = {data_out_rows[837*col_length-1 -: col_length]};
assign pixels_col_23_9 = {data_out_cols[838*col_length-1 -: col_length]};
assign pixels_row_23_9 = {data_out_rows[838*col_length-1 -: col_length]};
assign pixels_col_23_10 = {data_out_cols[839*col_length-1 -: col_length]};
assign pixels_row_23_10 = {data_out_rows[839*col_length-1 -: col_length]};
assign pixels_col_23_11 = {data_out_cols[840*col_length-1 -: col_length]};
assign pixels_row_23_11 = {data_out_rows[840*col_length-1 -: col_length]};
assign pixels_col_23_12 = {data_out_cols[841*col_length-1 -: col_length]};
assign pixels_row_23_12 = {data_out_rows[841*col_length-1 -: col_length]};
assign pixels_col_23_13 = {data_out_cols[842*col_length-1 -: col_length]};
assign pixels_row_23_13 = {data_out_rows[842*col_length-1 -: col_length]};
assign pixels_col_23_14 = {data_out_cols[843*col_length-1 -: col_length]};
assign pixels_row_23_14 = {data_out_rows[843*col_length-1 -: col_length]};
assign pixels_col_23_15 = {data_out_cols[844*col_length-1 -: col_length]};
assign pixels_row_23_15 = {data_out_rows[844*col_length-1 -: col_length]};
assign pixels_col_23_16 = {data_out_cols[845*col_length-1 -: col_length]};
assign pixels_row_23_16 = {data_out_rows[845*col_length-1 -: col_length]};
assign pixels_col_23_17 = {data_out_cols[846*col_length-1 -: col_length]};
assign pixels_row_23_17 = {data_out_rows[846*col_length-1 -: col_length]};
assign pixels_col_23_18 = {data_out_cols[847*col_length-1 -: col_length]};
assign pixels_row_23_18 = {data_out_rows[847*col_length-1 -: col_length]};
assign pixels_col_23_19 = {data_out_cols[848*col_length-1 -: col_length]};
assign pixels_row_23_19 = {data_out_rows[848*col_length-1 -: col_length]};
assign pixels_col_23_20 = {data_out_cols[849*col_length-1 -: col_length]};
assign pixels_row_23_20 = {data_out_rows[849*col_length-1 -: col_length]};
assign pixels_col_23_21 = {data_out_cols[850*col_length-1 -: col_length]};
assign pixels_row_23_21 = {data_out_rows[850*col_length-1 -: col_length]};
assign pixels_col_23_22 = {data_out_cols[851*col_length-1 -: col_length]};
assign pixels_row_23_22 = {data_out_rows[851*col_length-1 -: col_length]};
assign pixels_col_23_23 = {data_out_cols[852*col_length-1 -: col_length]};
assign pixels_row_23_23 = {data_out_rows[852*col_length-1 -: col_length]};
assign pixels_col_23_24 = {data_out_cols[853*col_length-1 -: col_length]};
assign pixels_row_23_24 = {data_out_rows[853*col_length-1 -: col_length]};
assign pixels_col_23_25 = {data_out_cols[854*col_length-1 -: col_length]};
assign pixels_row_23_25 = {data_out_rows[854*col_length-1 -: col_length]};
assign pixels_col_23_26 = {data_out_cols[855*col_length-1 -: col_length]};
assign pixels_row_23_26 = {data_out_rows[855*col_length-1 -: col_length]};
assign pixels_col_23_27 = {data_out_cols[856*col_length-1 -: col_length]};
assign pixels_row_23_27 = {data_out_rows[856*col_length-1 -: col_length]};
assign pixels_col_23_28 = {data_out_cols[857*col_length-1 -: col_length]};
assign pixels_row_23_28 = {data_out_rows[857*col_length-1 -: col_length]};
assign pixels_col_23_29 = {data_out_cols[858*col_length-1 -: col_length]};
assign pixels_row_23_29 = {data_out_rows[858*col_length-1 -: col_length]};
assign pixels_col_23_30 = {data_out_cols[859*col_length-1 -: col_length]};
assign pixels_row_23_30 = {data_out_rows[859*col_length-1 -: col_length]};
assign pixels_col_23_31 = {data_out_cols[860*col_length-1 -: col_length]};
assign pixels_row_23_31 = {data_out_rows[860*col_length-1 -: col_length]};
assign pixels_col_23_32 = {data_out_cols[861*col_length-1 -: col_length]};
assign pixels_row_23_32 = {data_out_rows[861*col_length-1 -: col_length]};
assign pixels_col_23_33 = {data_out_cols[862*col_length-1 -: col_length]};
assign pixels_row_23_33 = {data_out_rows[862*col_length-1 -: col_length]};
assign pixels_col_23_34 = {data_out_cols[863*col_length-1 -: col_length]};
assign pixels_row_23_34 = {data_out_rows[863*col_length-1 -: col_length]};
assign pixels_col_23_35 = {data_out_cols[864*col_length-1 -: col_length]};
assign pixels_row_23_35 = {data_out_rows[864*col_length-1 -: col_length]};
assign pixels_col_24_0 = {data_out_cols[865*col_length-1 -: col_length]};
assign pixels_row_24_0 = {data_out_rows[865*col_length-1 -: col_length]};
assign pixels_col_24_1 = {data_out_cols[866*col_length-1 -: col_length]};
assign pixels_row_24_1 = {data_out_rows[866*col_length-1 -: col_length]};
assign pixels_col_24_2 = {data_out_cols[867*col_length-1 -: col_length]};
assign pixels_row_24_2 = {data_out_rows[867*col_length-1 -: col_length]};
assign pixels_col_24_3 = {data_out_cols[868*col_length-1 -: col_length]};
assign pixels_row_24_3 = {data_out_rows[868*col_length-1 -: col_length]};
assign pixels_col_24_4 = {data_out_cols[869*col_length-1 -: col_length]};
assign pixels_row_24_4 = {data_out_rows[869*col_length-1 -: col_length]};
assign pixels_col_24_5 = {data_out_cols[870*col_length-1 -: col_length]};
assign pixels_row_24_5 = {data_out_rows[870*col_length-1 -: col_length]};
assign pixels_col_24_6 = {data_out_cols[871*col_length-1 -: col_length]};
assign pixels_row_24_6 = {data_out_rows[871*col_length-1 -: col_length]};
assign pixels_col_24_7 = {data_out_cols[872*col_length-1 -: col_length]};
assign pixels_row_24_7 = {data_out_rows[872*col_length-1 -: col_length]};
assign pixels_col_24_8 = {data_out_cols[873*col_length-1 -: col_length]};
assign pixels_row_24_8 = {data_out_rows[873*col_length-1 -: col_length]};
assign pixels_col_24_9 = {data_out_cols[874*col_length-1 -: col_length]};
assign pixels_row_24_9 = {data_out_rows[874*col_length-1 -: col_length]};
assign pixels_col_24_10 = {data_out_cols[875*col_length-1 -: col_length]};
assign pixels_row_24_10 = {data_out_rows[875*col_length-1 -: col_length]};
assign pixels_col_24_11 = {data_out_cols[876*col_length-1 -: col_length]};
assign pixels_row_24_11 = {data_out_rows[876*col_length-1 -: col_length]};
assign pixels_col_24_12 = {data_out_cols[877*col_length-1 -: col_length]};
assign pixels_row_24_12 = {data_out_rows[877*col_length-1 -: col_length]};
assign pixels_col_24_13 = {data_out_cols[878*col_length-1 -: col_length]};
assign pixels_row_24_13 = {data_out_rows[878*col_length-1 -: col_length]};
assign pixels_col_24_14 = {data_out_cols[879*col_length-1 -: col_length]};
assign pixels_row_24_14 = {data_out_rows[879*col_length-1 -: col_length]};
assign pixels_col_24_15 = {data_out_cols[880*col_length-1 -: col_length]};
assign pixels_row_24_15 = {data_out_rows[880*col_length-1 -: col_length]};
assign pixels_col_24_16 = {data_out_cols[881*col_length-1 -: col_length]};
assign pixels_row_24_16 = {data_out_rows[881*col_length-1 -: col_length]};
assign pixels_col_24_17 = {data_out_cols[882*col_length-1 -: col_length]};
assign pixels_row_24_17 = {data_out_rows[882*col_length-1 -: col_length]};
assign pixels_col_24_18 = {data_out_cols[883*col_length-1 -: col_length]};
assign pixels_row_24_18 = {data_out_rows[883*col_length-1 -: col_length]};
assign pixels_col_24_19 = {data_out_cols[884*col_length-1 -: col_length]};
assign pixels_row_24_19 = {data_out_rows[884*col_length-1 -: col_length]};
assign pixels_col_24_20 = {data_out_cols[885*col_length-1 -: col_length]};
assign pixels_row_24_20 = {data_out_rows[885*col_length-1 -: col_length]};
assign pixels_col_24_21 = {data_out_cols[886*col_length-1 -: col_length]};
assign pixels_row_24_21 = {data_out_rows[886*col_length-1 -: col_length]};
assign pixels_col_24_22 = {data_out_cols[887*col_length-1 -: col_length]};
assign pixels_row_24_22 = {data_out_rows[887*col_length-1 -: col_length]};
assign pixels_col_24_23 = {data_out_cols[888*col_length-1 -: col_length]};
assign pixels_row_24_23 = {data_out_rows[888*col_length-1 -: col_length]};
assign pixels_col_24_24 = {data_out_cols[889*col_length-1 -: col_length]};
assign pixels_row_24_24 = {data_out_rows[889*col_length-1 -: col_length]};
assign pixels_col_24_25 = {data_out_cols[890*col_length-1 -: col_length]};
assign pixels_row_24_25 = {data_out_rows[890*col_length-1 -: col_length]};
assign pixels_col_24_26 = {data_out_cols[891*col_length-1 -: col_length]};
assign pixels_row_24_26 = {data_out_rows[891*col_length-1 -: col_length]};
assign pixels_col_24_27 = {data_out_cols[892*col_length-1 -: col_length]};
assign pixels_row_24_27 = {data_out_rows[892*col_length-1 -: col_length]};
assign pixels_col_24_28 = {data_out_cols[893*col_length-1 -: col_length]};
assign pixels_row_24_28 = {data_out_rows[893*col_length-1 -: col_length]};
assign pixels_col_24_29 = {data_out_cols[894*col_length-1 -: col_length]};
assign pixels_row_24_29 = {data_out_rows[894*col_length-1 -: col_length]};
assign pixels_col_24_30 = {data_out_cols[895*col_length-1 -: col_length]};
assign pixels_row_24_30 = {data_out_rows[895*col_length-1 -: col_length]};
assign pixels_col_24_31 = {data_out_cols[896*col_length-1 -: col_length]};
assign pixels_row_24_31 = {data_out_rows[896*col_length-1 -: col_length]};
assign pixels_col_24_32 = {data_out_cols[897*col_length-1 -: col_length]};
assign pixels_row_24_32 = {data_out_rows[897*col_length-1 -: col_length]};
assign pixels_col_24_33 = {data_out_cols[898*col_length-1 -: col_length]};
assign pixels_row_24_33 = {data_out_rows[898*col_length-1 -: col_length]};
assign pixels_col_24_34 = {data_out_cols[899*col_length-1 -: col_length]};
assign pixels_row_24_34 = {data_out_rows[899*col_length-1 -: col_length]};
assign pixels_col_24_35 = {data_out_cols[900*col_length-1 -: col_length]};
assign pixels_row_24_35 = {data_out_rows[900*col_length-1 -: col_length]};
assign pixels_col_25_0 = {data_out_cols[901*col_length-1 -: col_length]};
assign pixels_row_25_0 = {data_out_rows[901*col_length-1 -: col_length]};
assign pixels_col_25_1 = {data_out_cols[902*col_length-1 -: col_length]};
assign pixels_row_25_1 = {data_out_rows[902*col_length-1 -: col_length]};
assign pixels_col_25_2 = {data_out_cols[903*col_length-1 -: col_length]};
assign pixels_row_25_2 = {data_out_rows[903*col_length-1 -: col_length]};
assign pixels_col_25_3 = {data_out_cols[904*col_length-1 -: col_length]};
assign pixels_row_25_3 = {data_out_rows[904*col_length-1 -: col_length]};
assign pixels_col_25_4 = {data_out_cols[905*col_length-1 -: col_length]};
assign pixels_row_25_4 = {data_out_rows[905*col_length-1 -: col_length]};
assign pixels_col_25_5 = {data_out_cols[906*col_length-1 -: col_length]};
assign pixels_row_25_5 = {data_out_rows[906*col_length-1 -: col_length]};
assign pixels_col_25_6 = {data_out_cols[907*col_length-1 -: col_length]};
assign pixels_row_25_6 = {data_out_rows[907*col_length-1 -: col_length]};
assign pixels_col_25_7 = {data_out_cols[908*col_length-1 -: col_length]};
assign pixels_row_25_7 = {data_out_rows[908*col_length-1 -: col_length]};
assign pixels_col_25_8 = {data_out_cols[909*col_length-1 -: col_length]};
assign pixels_row_25_8 = {data_out_rows[909*col_length-1 -: col_length]};
assign pixels_col_25_9 = {data_out_cols[910*col_length-1 -: col_length]};
assign pixels_row_25_9 = {data_out_rows[910*col_length-1 -: col_length]};
assign pixels_col_25_10 = {data_out_cols[911*col_length-1 -: col_length]};
assign pixels_row_25_10 = {data_out_rows[911*col_length-1 -: col_length]};
assign pixels_col_25_11 = {data_out_cols[912*col_length-1 -: col_length]};
assign pixels_row_25_11 = {data_out_rows[912*col_length-1 -: col_length]};
assign pixels_col_25_12 = {data_out_cols[913*col_length-1 -: col_length]};
assign pixels_row_25_12 = {data_out_rows[913*col_length-1 -: col_length]};
assign pixels_col_25_13 = {data_out_cols[914*col_length-1 -: col_length]};
assign pixels_row_25_13 = {data_out_rows[914*col_length-1 -: col_length]};
assign pixels_col_25_14 = {data_out_cols[915*col_length-1 -: col_length]};
assign pixels_row_25_14 = {data_out_rows[915*col_length-1 -: col_length]};
assign pixels_col_25_15 = {data_out_cols[916*col_length-1 -: col_length]};
assign pixels_row_25_15 = {data_out_rows[916*col_length-1 -: col_length]};
assign pixels_col_25_16 = {data_out_cols[917*col_length-1 -: col_length]};
assign pixels_row_25_16 = {data_out_rows[917*col_length-1 -: col_length]};
assign pixels_col_25_17 = {data_out_cols[918*col_length-1 -: col_length]};
assign pixels_row_25_17 = {data_out_rows[918*col_length-1 -: col_length]};
assign pixels_col_25_18 = {data_out_cols[919*col_length-1 -: col_length]};
assign pixels_row_25_18 = {data_out_rows[919*col_length-1 -: col_length]};
assign pixels_col_25_19 = {data_out_cols[920*col_length-1 -: col_length]};
assign pixels_row_25_19 = {data_out_rows[920*col_length-1 -: col_length]};
assign pixels_col_25_20 = {data_out_cols[921*col_length-1 -: col_length]};
assign pixels_row_25_20 = {data_out_rows[921*col_length-1 -: col_length]};
assign pixels_col_25_21 = {data_out_cols[922*col_length-1 -: col_length]};
assign pixels_row_25_21 = {data_out_rows[922*col_length-1 -: col_length]};
assign pixels_col_25_22 = {data_out_cols[923*col_length-1 -: col_length]};
assign pixels_row_25_22 = {data_out_rows[923*col_length-1 -: col_length]};
assign pixels_col_25_23 = {data_out_cols[924*col_length-1 -: col_length]};
assign pixels_row_25_23 = {data_out_rows[924*col_length-1 -: col_length]};
assign pixels_col_25_24 = {data_out_cols[925*col_length-1 -: col_length]};
assign pixels_row_25_24 = {data_out_rows[925*col_length-1 -: col_length]};
assign pixels_col_25_25 = {data_out_cols[926*col_length-1 -: col_length]};
assign pixels_row_25_25 = {data_out_rows[926*col_length-1 -: col_length]};
assign pixels_col_25_26 = {data_out_cols[927*col_length-1 -: col_length]};
assign pixels_row_25_26 = {data_out_rows[927*col_length-1 -: col_length]};
assign pixels_col_25_27 = {data_out_cols[928*col_length-1 -: col_length]};
assign pixels_row_25_27 = {data_out_rows[928*col_length-1 -: col_length]};
assign pixels_col_25_28 = {data_out_cols[929*col_length-1 -: col_length]};
assign pixels_row_25_28 = {data_out_rows[929*col_length-1 -: col_length]};
assign pixels_col_25_29 = {data_out_cols[930*col_length-1 -: col_length]};
assign pixels_row_25_29 = {data_out_rows[930*col_length-1 -: col_length]};
assign pixels_col_25_30 = {data_out_cols[931*col_length-1 -: col_length]};
assign pixels_row_25_30 = {data_out_rows[931*col_length-1 -: col_length]};
assign pixels_col_25_31 = {data_out_cols[932*col_length-1 -: col_length]};
assign pixels_row_25_31 = {data_out_rows[932*col_length-1 -: col_length]};
assign pixels_col_25_32 = {data_out_cols[933*col_length-1 -: col_length]};
assign pixels_row_25_32 = {data_out_rows[933*col_length-1 -: col_length]};
assign pixels_col_25_33 = {data_out_cols[934*col_length-1 -: col_length]};
assign pixels_row_25_33 = {data_out_rows[934*col_length-1 -: col_length]};
assign pixels_col_25_34 = {data_out_cols[935*col_length-1 -: col_length]};
assign pixels_row_25_34 = {data_out_rows[935*col_length-1 -: col_length]};
assign pixels_col_25_35 = {data_out_cols[936*col_length-1 -: col_length]};
assign pixels_row_25_35 = {data_out_rows[936*col_length-1 -: col_length]};
assign pixels_col_26_0 = {data_out_cols[937*col_length-1 -: col_length]};
assign pixels_row_26_0 = {data_out_rows[937*col_length-1 -: col_length]};
assign pixels_col_26_1 = {data_out_cols[938*col_length-1 -: col_length]};
assign pixels_row_26_1 = {data_out_rows[938*col_length-1 -: col_length]};
assign pixels_col_26_2 = {data_out_cols[939*col_length-1 -: col_length]};
assign pixels_row_26_2 = {data_out_rows[939*col_length-1 -: col_length]};
assign pixels_col_26_3 = {data_out_cols[940*col_length-1 -: col_length]};
assign pixels_row_26_3 = {data_out_rows[940*col_length-1 -: col_length]};
assign pixels_col_26_4 = {data_out_cols[941*col_length-1 -: col_length]};
assign pixels_row_26_4 = {data_out_rows[941*col_length-1 -: col_length]};
assign pixels_col_26_5 = {data_out_cols[942*col_length-1 -: col_length]};
assign pixels_row_26_5 = {data_out_rows[942*col_length-1 -: col_length]};
assign pixels_col_26_6 = {data_out_cols[943*col_length-1 -: col_length]};
assign pixels_row_26_6 = {data_out_rows[943*col_length-1 -: col_length]};
assign pixels_col_26_7 = {data_out_cols[944*col_length-1 -: col_length]};
assign pixels_row_26_7 = {data_out_rows[944*col_length-1 -: col_length]};
assign pixels_col_26_8 = {data_out_cols[945*col_length-1 -: col_length]};
assign pixels_row_26_8 = {data_out_rows[945*col_length-1 -: col_length]};
assign pixels_col_26_9 = {data_out_cols[946*col_length-1 -: col_length]};
assign pixels_row_26_9 = {data_out_rows[946*col_length-1 -: col_length]};
assign pixels_col_26_10 = {data_out_cols[947*col_length-1 -: col_length]};
assign pixels_row_26_10 = {data_out_rows[947*col_length-1 -: col_length]};
assign pixels_col_26_11 = {data_out_cols[948*col_length-1 -: col_length]};
assign pixels_row_26_11 = {data_out_rows[948*col_length-1 -: col_length]};
assign pixels_col_26_12 = {data_out_cols[949*col_length-1 -: col_length]};
assign pixels_row_26_12 = {data_out_rows[949*col_length-1 -: col_length]};
assign pixels_col_26_13 = {data_out_cols[950*col_length-1 -: col_length]};
assign pixels_row_26_13 = {data_out_rows[950*col_length-1 -: col_length]};
assign pixels_col_26_14 = {data_out_cols[951*col_length-1 -: col_length]};
assign pixels_row_26_14 = {data_out_rows[951*col_length-1 -: col_length]};
assign pixels_col_26_15 = {data_out_cols[952*col_length-1 -: col_length]};
assign pixels_row_26_15 = {data_out_rows[952*col_length-1 -: col_length]};
assign pixels_col_26_16 = {data_out_cols[953*col_length-1 -: col_length]};
assign pixels_row_26_16 = {data_out_rows[953*col_length-1 -: col_length]};
assign pixels_col_26_17 = {data_out_cols[954*col_length-1 -: col_length]};
assign pixels_row_26_17 = {data_out_rows[954*col_length-1 -: col_length]};
assign pixels_col_26_18 = {data_out_cols[955*col_length-1 -: col_length]};
assign pixels_row_26_18 = {data_out_rows[955*col_length-1 -: col_length]};
assign pixels_col_26_19 = {data_out_cols[956*col_length-1 -: col_length]};
assign pixels_row_26_19 = {data_out_rows[956*col_length-1 -: col_length]};
assign pixels_col_26_20 = {data_out_cols[957*col_length-1 -: col_length]};
assign pixels_row_26_20 = {data_out_rows[957*col_length-1 -: col_length]};
assign pixels_col_26_21 = {data_out_cols[958*col_length-1 -: col_length]};
assign pixels_row_26_21 = {data_out_rows[958*col_length-1 -: col_length]};
assign pixels_col_26_22 = {data_out_cols[959*col_length-1 -: col_length]};
assign pixels_row_26_22 = {data_out_rows[959*col_length-1 -: col_length]};
assign pixels_col_26_23 = {data_out_cols[960*col_length-1 -: col_length]};
assign pixels_row_26_23 = {data_out_rows[960*col_length-1 -: col_length]};
assign pixels_col_26_24 = {data_out_cols[961*col_length-1 -: col_length]};
assign pixels_row_26_24 = {data_out_rows[961*col_length-1 -: col_length]};
assign pixels_col_26_25 = {data_out_cols[962*col_length-1 -: col_length]};
assign pixels_row_26_25 = {data_out_rows[962*col_length-1 -: col_length]};
assign pixels_col_26_26 = {data_out_cols[963*col_length-1 -: col_length]};
assign pixels_row_26_26 = {data_out_rows[963*col_length-1 -: col_length]};
assign pixels_col_26_27 = {data_out_cols[964*col_length-1 -: col_length]};
assign pixels_row_26_27 = {data_out_rows[964*col_length-1 -: col_length]};
assign pixels_col_26_28 = {data_out_cols[965*col_length-1 -: col_length]};
assign pixels_row_26_28 = {data_out_rows[965*col_length-1 -: col_length]};
assign pixels_col_26_29 = {data_out_cols[966*col_length-1 -: col_length]};
assign pixels_row_26_29 = {data_out_rows[966*col_length-1 -: col_length]};
assign pixels_col_26_30 = {data_out_cols[967*col_length-1 -: col_length]};
assign pixels_row_26_30 = {data_out_rows[967*col_length-1 -: col_length]};
assign pixels_col_26_31 = {data_out_cols[968*col_length-1 -: col_length]};
assign pixels_row_26_31 = {data_out_rows[968*col_length-1 -: col_length]};
assign pixels_col_26_32 = {data_out_cols[969*col_length-1 -: col_length]};
assign pixels_row_26_32 = {data_out_rows[969*col_length-1 -: col_length]};
assign pixels_col_26_33 = {data_out_cols[970*col_length-1 -: col_length]};
assign pixels_row_26_33 = {data_out_rows[970*col_length-1 -: col_length]};
assign pixels_col_26_34 = {data_out_cols[971*col_length-1 -: col_length]};
assign pixels_row_26_34 = {data_out_rows[971*col_length-1 -: col_length]};
assign pixels_col_26_35 = {data_out_cols[972*col_length-1 -: col_length]};
assign pixels_row_26_35 = {data_out_rows[972*col_length-1 -: col_length]};
assign pixels_col_27_0 = {data_out_cols[973*col_length-1 -: col_length]};
assign pixels_row_27_0 = {data_out_rows[973*col_length-1 -: col_length]};
assign pixels_col_27_1 = {data_out_cols[974*col_length-1 -: col_length]};
assign pixels_row_27_1 = {data_out_rows[974*col_length-1 -: col_length]};
assign pixels_col_27_2 = {data_out_cols[975*col_length-1 -: col_length]};
assign pixels_row_27_2 = {data_out_rows[975*col_length-1 -: col_length]};
assign pixels_col_27_3 = {data_out_cols[976*col_length-1 -: col_length]};
assign pixels_row_27_3 = {data_out_rows[976*col_length-1 -: col_length]};
assign pixels_col_27_4 = {data_out_cols[977*col_length-1 -: col_length]};
assign pixels_row_27_4 = {data_out_rows[977*col_length-1 -: col_length]};
assign pixels_col_27_5 = {data_out_cols[978*col_length-1 -: col_length]};
assign pixels_row_27_5 = {data_out_rows[978*col_length-1 -: col_length]};
assign pixels_col_27_6 = {data_out_cols[979*col_length-1 -: col_length]};
assign pixels_row_27_6 = {data_out_rows[979*col_length-1 -: col_length]};
assign pixels_col_27_7 = {data_out_cols[980*col_length-1 -: col_length]};
assign pixels_row_27_7 = {data_out_rows[980*col_length-1 -: col_length]};
assign pixels_col_27_8 = {data_out_cols[981*col_length-1 -: col_length]};
assign pixels_row_27_8 = {data_out_rows[981*col_length-1 -: col_length]};
assign pixels_col_27_9 = {data_out_cols[982*col_length-1 -: col_length]};
assign pixels_row_27_9 = {data_out_rows[982*col_length-1 -: col_length]};
assign pixels_col_27_10 = {data_out_cols[983*col_length-1 -: col_length]};
assign pixels_row_27_10 = {data_out_rows[983*col_length-1 -: col_length]};
assign pixels_col_27_11 = {data_out_cols[984*col_length-1 -: col_length]};
assign pixels_row_27_11 = {data_out_rows[984*col_length-1 -: col_length]};
assign pixels_col_27_12 = {data_out_cols[985*col_length-1 -: col_length]};
assign pixels_row_27_12 = {data_out_rows[985*col_length-1 -: col_length]};
assign pixels_col_27_13 = {data_out_cols[986*col_length-1 -: col_length]};
assign pixels_row_27_13 = {data_out_rows[986*col_length-1 -: col_length]};
assign pixels_col_27_14 = {data_out_cols[987*col_length-1 -: col_length]};
assign pixels_row_27_14 = {data_out_rows[987*col_length-1 -: col_length]};
assign pixels_col_27_15 = {data_out_cols[988*col_length-1 -: col_length]};
assign pixels_row_27_15 = {data_out_rows[988*col_length-1 -: col_length]};
assign pixels_col_27_16 = {data_out_cols[989*col_length-1 -: col_length]};
assign pixels_row_27_16 = {data_out_rows[989*col_length-1 -: col_length]};
assign pixels_col_27_17 = {data_out_cols[990*col_length-1 -: col_length]};
assign pixels_row_27_17 = {data_out_rows[990*col_length-1 -: col_length]};
assign pixels_col_27_18 = {data_out_cols[991*col_length-1 -: col_length]};
assign pixels_row_27_18 = {data_out_rows[991*col_length-1 -: col_length]};
assign pixels_col_27_19 = {data_out_cols[992*col_length-1 -: col_length]};
assign pixels_row_27_19 = {data_out_rows[992*col_length-1 -: col_length]};
assign pixels_col_27_20 = {data_out_cols[993*col_length-1 -: col_length]};
assign pixels_row_27_20 = {data_out_rows[993*col_length-1 -: col_length]};
assign pixels_col_27_21 = {data_out_cols[994*col_length-1 -: col_length]};
assign pixels_row_27_21 = {data_out_rows[994*col_length-1 -: col_length]};
assign pixels_col_27_22 = {data_out_cols[995*col_length-1 -: col_length]};
assign pixels_row_27_22 = {data_out_rows[995*col_length-1 -: col_length]};
assign pixels_col_27_23 = {data_out_cols[996*col_length-1 -: col_length]};
assign pixels_row_27_23 = {data_out_rows[996*col_length-1 -: col_length]};
assign pixels_col_27_24 = {data_out_cols[997*col_length-1 -: col_length]};
assign pixels_row_27_24 = {data_out_rows[997*col_length-1 -: col_length]};
assign pixels_col_27_25 = {data_out_cols[998*col_length-1 -: col_length]};
assign pixels_row_27_25 = {data_out_rows[998*col_length-1 -: col_length]};
assign pixels_col_27_26 = {data_out_cols[999*col_length-1 -: col_length]};
assign pixels_row_27_26 = {data_out_rows[999*col_length-1 -: col_length]};
assign pixels_col_27_27 = {data_out_cols[1000*col_length-1 -: col_length]};
assign pixels_row_27_27 = {data_out_rows[1000*col_length-1 -: col_length]};
assign pixels_col_27_28 = {data_out_cols[1001*col_length-1 -: col_length]};
assign pixels_row_27_28 = {data_out_rows[1001*col_length-1 -: col_length]};
assign pixels_col_27_29 = {data_out_cols[1002*col_length-1 -: col_length]};
assign pixels_row_27_29 = {data_out_rows[1002*col_length-1 -: col_length]};
assign pixels_col_27_30 = {data_out_cols[1003*col_length-1 -: col_length]};
assign pixels_row_27_30 = {data_out_rows[1003*col_length-1 -: col_length]};
assign pixels_col_27_31 = {data_out_cols[1004*col_length-1 -: col_length]};
assign pixels_row_27_31 = {data_out_rows[1004*col_length-1 -: col_length]};
assign pixels_col_27_32 = {data_out_cols[1005*col_length-1 -: col_length]};
assign pixels_row_27_32 = {data_out_rows[1005*col_length-1 -: col_length]};
assign pixels_col_27_33 = {data_out_cols[1006*col_length-1 -: col_length]};
assign pixels_row_27_33 = {data_out_rows[1006*col_length-1 -: col_length]};
assign pixels_col_27_34 = {data_out_cols[1007*col_length-1 -: col_length]};
assign pixels_row_27_34 = {data_out_rows[1007*col_length-1 -: col_length]};
assign pixels_col_27_35 = {data_out_cols[1008*col_length-1 -: col_length]};
assign pixels_row_27_35 = {data_out_rows[1008*col_length-1 -: col_length]};
assign pixels_col_28_0 = {data_out_cols[1009*col_length-1 -: col_length]};
assign pixels_row_28_0 = {data_out_rows[1009*col_length-1 -: col_length]};
assign pixels_col_28_1 = {data_out_cols[1010*col_length-1 -: col_length]};
assign pixels_row_28_1 = {data_out_rows[1010*col_length-1 -: col_length]};
assign pixels_col_28_2 = {data_out_cols[1011*col_length-1 -: col_length]};
assign pixels_row_28_2 = {data_out_rows[1011*col_length-1 -: col_length]};
assign pixels_col_28_3 = {data_out_cols[1012*col_length-1 -: col_length]};
assign pixels_row_28_3 = {data_out_rows[1012*col_length-1 -: col_length]};
assign pixels_col_28_4 = {data_out_cols[1013*col_length-1 -: col_length]};
assign pixels_row_28_4 = {data_out_rows[1013*col_length-1 -: col_length]};
assign pixels_col_28_5 = {data_out_cols[1014*col_length-1 -: col_length]};
assign pixels_row_28_5 = {data_out_rows[1014*col_length-1 -: col_length]};
assign pixels_col_28_6 = {data_out_cols[1015*col_length-1 -: col_length]};
assign pixels_row_28_6 = {data_out_rows[1015*col_length-1 -: col_length]};
assign pixels_col_28_7 = {data_out_cols[1016*col_length-1 -: col_length]};
assign pixels_row_28_7 = {data_out_rows[1016*col_length-1 -: col_length]};
assign pixels_col_28_8 = {data_out_cols[1017*col_length-1 -: col_length]};
assign pixels_row_28_8 = {data_out_rows[1017*col_length-1 -: col_length]};
assign pixels_col_28_9 = {data_out_cols[1018*col_length-1 -: col_length]};
assign pixels_row_28_9 = {data_out_rows[1018*col_length-1 -: col_length]};
assign pixels_col_28_10 = {data_out_cols[1019*col_length-1 -: col_length]};
assign pixels_row_28_10 = {data_out_rows[1019*col_length-1 -: col_length]};
assign pixels_col_28_11 = {data_out_cols[1020*col_length-1 -: col_length]};
assign pixels_row_28_11 = {data_out_rows[1020*col_length-1 -: col_length]};
assign pixels_col_28_12 = {data_out_cols[1021*col_length-1 -: col_length]};
assign pixels_row_28_12 = {data_out_rows[1021*col_length-1 -: col_length]};
assign pixels_col_28_13 = {data_out_cols[1022*col_length-1 -: col_length]};
assign pixels_row_28_13 = {data_out_rows[1022*col_length-1 -: col_length]};
assign pixels_col_28_14 = {data_out_cols[1023*col_length-1 -: col_length]};
assign pixels_row_28_14 = {data_out_rows[1023*col_length-1 -: col_length]};
assign pixels_col_28_15 = {data_out_cols[1024*col_length-1 -: col_length]};
assign pixels_row_28_15 = {data_out_rows[1024*col_length-1 -: col_length]};
assign pixels_col_28_16 = {data_out_cols[1025*col_length-1 -: col_length]};
assign pixels_row_28_16 = {data_out_rows[1025*col_length-1 -: col_length]};
assign pixels_col_28_17 = {data_out_cols[1026*col_length-1 -: col_length]};
assign pixels_row_28_17 = {data_out_rows[1026*col_length-1 -: col_length]};
assign pixels_col_28_18 = {data_out_cols[1027*col_length-1 -: col_length]};
assign pixels_row_28_18 = {data_out_rows[1027*col_length-1 -: col_length]};
assign pixels_col_28_19 = {data_out_cols[1028*col_length-1 -: col_length]};
assign pixels_row_28_19 = {data_out_rows[1028*col_length-1 -: col_length]};
assign pixels_col_28_20 = {data_out_cols[1029*col_length-1 -: col_length]};
assign pixels_row_28_20 = {data_out_rows[1029*col_length-1 -: col_length]};
assign pixels_col_28_21 = {data_out_cols[1030*col_length-1 -: col_length]};
assign pixels_row_28_21 = {data_out_rows[1030*col_length-1 -: col_length]};
assign pixels_col_28_22 = {data_out_cols[1031*col_length-1 -: col_length]};
assign pixels_row_28_22 = {data_out_rows[1031*col_length-1 -: col_length]};
assign pixels_col_28_23 = {data_out_cols[1032*col_length-1 -: col_length]};
assign pixels_row_28_23 = {data_out_rows[1032*col_length-1 -: col_length]};
assign pixels_col_28_24 = {data_out_cols[1033*col_length-1 -: col_length]};
assign pixels_row_28_24 = {data_out_rows[1033*col_length-1 -: col_length]};
assign pixels_col_28_25 = {data_out_cols[1034*col_length-1 -: col_length]};
assign pixels_row_28_25 = {data_out_rows[1034*col_length-1 -: col_length]};
assign pixels_col_28_26 = {data_out_cols[1035*col_length-1 -: col_length]};
assign pixels_row_28_26 = {data_out_rows[1035*col_length-1 -: col_length]};
assign pixels_col_28_27 = {data_out_cols[1036*col_length-1 -: col_length]};
assign pixels_row_28_27 = {data_out_rows[1036*col_length-1 -: col_length]};
assign pixels_col_28_28 = {data_out_cols[1037*col_length-1 -: col_length]};
assign pixels_row_28_28 = {data_out_rows[1037*col_length-1 -: col_length]};
assign pixels_col_28_29 = {data_out_cols[1038*col_length-1 -: col_length]};
assign pixels_row_28_29 = {data_out_rows[1038*col_length-1 -: col_length]};
assign pixels_col_28_30 = {data_out_cols[1039*col_length-1 -: col_length]};
assign pixels_row_28_30 = {data_out_rows[1039*col_length-1 -: col_length]};
assign pixels_col_28_31 = {data_out_cols[1040*col_length-1 -: col_length]};
assign pixels_row_28_31 = {data_out_rows[1040*col_length-1 -: col_length]};
assign pixels_col_28_32 = {data_out_cols[1041*col_length-1 -: col_length]};
assign pixels_row_28_32 = {data_out_rows[1041*col_length-1 -: col_length]};
assign pixels_col_28_33 = {data_out_cols[1042*col_length-1 -: col_length]};
assign pixels_row_28_33 = {data_out_rows[1042*col_length-1 -: col_length]};
assign pixels_col_28_34 = {data_out_cols[1043*col_length-1 -: col_length]};
assign pixels_row_28_34 = {data_out_rows[1043*col_length-1 -: col_length]};
assign pixels_col_28_35 = {data_out_cols[1044*col_length-1 -: col_length]};
assign pixels_row_28_35 = {data_out_rows[1044*col_length-1 -: col_length]};
assign pixels_col_29_0 = {data_out_cols[1045*col_length-1 -: col_length]};
assign pixels_row_29_0 = {data_out_rows[1045*col_length-1 -: col_length]};
assign pixels_col_29_1 = {data_out_cols[1046*col_length-1 -: col_length]};
assign pixels_row_29_1 = {data_out_rows[1046*col_length-1 -: col_length]};
assign pixels_col_29_2 = {data_out_cols[1047*col_length-1 -: col_length]};
assign pixels_row_29_2 = {data_out_rows[1047*col_length-1 -: col_length]};
assign pixels_col_29_3 = {data_out_cols[1048*col_length-1 -: col_length]};
assign pixels_row_29_3 = {data_out_rows[1048*col_length-1 -: col_length]};
assign pixels_col_29_4 = {data_out_cols[1049*col_length-1 -: col_length]};
assign pixels_row_29_4 = {data_out_rows[1049*col_length-1 -: col_length]};
assign pixels_col_29_5 = {data_out_cols[1050*col_length-1 -: col_length]};
assign pixels_row_29_5 = {data_out_rows[1050*col_length-1 -: col_length]};
assign pixels_col_29_6 = {data_out_cols[1051*col_length-1 -: col_length]};
assign pixels_row_29_6 = {data_out_rows[1051*col_length-1 -: col_length]};
assign pixels_col_29_7 = {data_out_cols[1052*col_length-1 -: col_length]};
assign pixels_row_29_7 = {data_out_rows[1052*col_length-1 -: col_length]};
assign pixels_col_29_8 = {data_out_cols[1053*col_length-1 -: col_length]};
assign pixels_row_29_8 = {data_out_rows[1053*col_length-1 -: col_length]};
assign pixels_col_29_9 = {data_out_cols[1054*col_length-1 -: col_length]};
assign pixels_row_29_9 = {data_out_rows[1054*col_length-1 -: col_length]};
assign pixels_col_29_10 = {data_out_cols[1055*col_length-1 -: col_length]};
assign pixels_row_29_10 = {data_out_rows[1055*col_length-1 -: col_length]};
assign pixels_col_29_11 = {data_out_cols[1056*col_length-1 -: col_length]};
assign pixels_row_29_11 = {data_out_rows[1056*col_length-1 -: col_length]};
assign pixels_col_29_12 = {data_out_cols[1057*col_length-1 -: col_length]};
assign pixels_row_29_12 = {data_out_rows[1057*col_length-1 -: col_length]};
assign pixels_col_29_13 = {data_out_cols[1058*col_length-1 -: col_length]};
assign pixels_row_29_13 = {data_out_rows[1058*col_length-1 -: col_length]};
assign pixels_col_29_14 = {data_out_cols[1059*col_length-1 -: col_length]};
assign pixels_row_29_14 = {data_out_rows[1059*col_length-1 -: col_length]};
assign pixels_col_29_15 = {data_out_cols[1060*col_length-1 -: col_length]};
assign pixels_row_29_15 = {data_out_rows[1060*col_length-1 -: col_length]};
assign pixels_col_29_16 = {data_out_cols[1061*col_length-1 -: col_length]};
assign pixels_row_29_16 = {data_out_rows[1061*col_length-1 -: col_length]};
assign pixels_col_29_17 = {data_out_cols[1062*col_length-1 -: col_length]};
assign pixels_row_29_17 = {data_out_rows[1062*col_length-1 -: col_length]};
assign pixels_col_29_18 = {data_out_cols[1063*col_length-1 -: col_length]};
assign pixels_row_29_18 = {data_out_rows[1063*col_length-1 -: col_length]};
assign pixels_col_29_19 = {data_out_cols[1064*col_length-1 -: col_length]};
assign pixels_row_29_19 = {data_out_rows[1064*col_length-1 -: col_length]};
assign pixels_col_29_20 = {data_out_cols[1065*col_length-1 -: col_length]};
assign pixels_row_29_20 = {data_out_rows[1065*col_length-1 -: col_length]};
assign pixels_col_29_21 = {data_out_cols[1066*col_length-1 -: col_length]};
assign pixels_row_29_21 = {data_out_rows[1066*col_length-1 -: col_length]};
assign pixels_col_29_22 = {data_out_cols[1067*col_length-1 -: col_length]};
assign pixels_row_29_22 = {data_out_rows[1067*col_length-1 -: col_length]};
assign pixels_col_29_23 = {data_out_cols[1068*col_length-1 -: col_length]};
assign pixels_row_29_23 = {data_out_rows[1068*col_length-1 -: col_length]};
assign pixels_col_29_24 = {data_out_cols[1069*col_length-1 -: col_length]};
assign pixels_row_29_24 = {data_out_rows[1069*col_length-1 -: col_length]};
assign pixels_col_29_25 = {data_out_cols[1070*col_length-1 -: col_length]};
assign pixels_row_29_25 = {data_out_rows[1070*col_length-1 -: col_length]};
assign pixels_col_29_26 = {data_out_cols[1071*col_length-1 -: col_length]};
assign pixels_row_29_26 = {data_out_rows[1071*col_length-1 -: col_length]};
assign pixels_col_29_27 = {data_out_cols[1072*col_length-1 -: col_length]};
assign pixels_row_29_27 = {data_out_rows[1072*col_length-1 -: col_length]};
assign pixels_col_29_28 = {data_out_cols[1073*col_length-1 -: col_length]};
assign pixels_row_29_28 = {data_out_rows[1073*col_length-1 -: col_length]};
assign pixels_col_29_29 = {data_out_cols[1074*col_length-1 -: col_length]};
assign pixels_row_29_29 = {data_out_rows[1074*col_length-1 -: col_length]};
assign pixels_col_29_30 = {data_out_cols[1075*col_length-1 -: col_length]};
assign pixels_row_29_30 = {data_out_rows[1075*col_length-1 -: col_length]};
assign pixels_col_29_31 = {data_out_cols[1076*col_length-1 -: col_length]};
assign pixels_row_29_31 = {data_out_rows[1076*col_length-1 -: col_length]};
assign pixels_col_29_32 = {data_out_cols[1077*col_length-1 -: col_length]};
assign pixels_row_29_32 = {data_out_rows[1077*col_length-1 -: col_length]};
assign pixels_col_29_33 = {data_out_cols[1078*col_length-1 -: col_length]};
assign pixels_row_29_33 = {data_out_rows[1078*col_length-1 -: col_length]};
assign pixels_col_29_34 = {data_out_cols[1079*col_length-1 -: col_length]};
assign pixels_row_29_34 = {data_out_rows[1079*col_length-1 -: col_length]};
assign pixels_col_29_35 = {data_out_cols[1080*col_length-1 -: col_length]};
assign pixels_row_29_35 = {data_out_rows[1080*col_length-1 -: col_length]};
assign pixels_col_30_0 = {data_out_cols[1081*col_length-1 -: col_length]};
assign pixels_row_30_0 = {data_out_rows[1081*col_length-1 -: col_length]};
assign pixels_col_30_1 = {data_out_cols[1082*col_length-1 -: col_length]};
assign pixels_row_30_1 = {data_out_rows[1082*col_length-1 -: col_length]};
assign pixels_col_30_2 = {data_out_cols[1083*col_length-1 -: col_length]};
assign pixels_row_30_2 = {data_out_rows[1083*col_length-1 -: col_length]};
assign pixels_col_30_3 = {data_out_cols[1084*col_length-1 -: col_length]};
assign pixels_row_30_3 = {data_out_rows[1084*col_length-1 -: col_length]};
assign pixels_col_30_4 = {data_out_cols[1085*col_length-1 -: col_length]};
assign pixels_row_30_4 = {data_out_rows[1085*col_length-1 -: col_length]};
assign pixels_col_30_5 = {data_out_cols[1086*col_length-1 -: col_length]};
assign pixels_row_30_5 = {data_out_rows[1086*col_length-1 -: col_length]};
assign pixels_col_30_6 = {data_out_cols[1087*col_length-1 -: col_length]};
assign pixels_row_30_6 = {data_out_rows[1087*col_length-1 -: col_length]};
assign pixels_col_30_7 = {data_out_cols[1088*col_length-1 -: col_length]};
assign pixels_row_30_7 = {data_out_rows[1088*col_length-1 -: col_length]};
assign pixels_col_30_8 = {data_out_cols[1089*col_length-1 -: col_length]};
assign pixels_row_30_8 = {data_out_rows[1089*col_length-1 -: col_length]};
assign pixels_col_30_9 = {data_out_cols[1090*col_length-1 -: col_length]};
assign pixels_row_30_9 = {data_out_rows[1090*col_length-1 -: col_length]};
assign pixels_col_30_10 = {data_out_cols[1091*col_length-1 -: col_length]};
assign pixels_row_30_10 = {data_out_rows[1091*col_length-1 -: col_length]};
assign pixels_col_30_11 = {data_out_cols[1092*col_length-1 -: col_length]};
assign pixels_row_30_11 = {data_out_rows[1092*col_length-1 -: col_length]};
assign pixels_col_30_12 = {data_out_cols[1093*col_length-1 -: col_length]};
assign pixels_row_30_12 = {data_out_rows[1093*col_length-1 -: col_length]};
assign pixels_col_30_13 = {data_out_cols[1094*col_length-1 -: col_length]};
assign pixels_row_30_13 = {data_out_rows[1094*col_length-1 -: col_length]};
assign pixels_col_30_14 = {data_out_cols[1095*col_length-1 -: col_length]};
assign pixels_row_30_14 = {data_out_rows[1095*col_length-1 -: col_length]};
assign pixels_col_30_15 = {data_out_cols[1096*col_length-1 -: col_length]};
assign pixels_row_30_15 = {data_out_rows[1096*col_length-1 -: col_length]};
assign pixels_col_30_16 = {data_out_cols[1097*col_length-1 -: col_length]};
assign pixels_row_30_16 = {data_out_rows[1097*col_length-1 -: col_length]};
assign pixels_col_30_17 = {data_out_cols[1098*col_length-1 -: col_length]};
assign pixels_row_30_17 = {data_out_rows[1098*col_length-1 -: col_length]};
assign pixels_col_30_18 = {data_out_cols[1099*col_length-1 -: col_length]};
assign pixels_row_30_18 = {data_out_rows[1099*col_length-1 -: col_length]};
assign pixels_col_30_19 = {data_out_cols[1100*col_length-1 -: col_length]};
assign pixels_row_30_19 = {data_out_rows[1100*col_length-1 -: col_length]};
assign pixels_col_30_20 = {data_out_cols[1101*col_length-1 -: col_length]};
assign pixels_row_30_20 = {data_out_rows[1101*col_length-1 -: col_length]};
assign pixels_col_30_21 = {data_out_cols[1102*col_length-1 -: col_length]};
assign pixels_row_30_21 = {data_out_rows[1102*col_length-1 -: col_length]};
assign pixels_col_30_22 = {data_out_cols[1103*col_length-1 -: col_length]};
assign pixels_row_30_22 = {data_out_rows[1103*col_length-1 -: col_length]};
assign pixels_col_30_23 = {data_out_cols[1104*col_length-1 -: col_length]};
assign pixels_row_30_23 = {data_out_rows[1104*col_length-1 -: col_length]};
assign pixels_col_30_24 = {data_out_cols[1105*col_length-1 -: col_length]};
assign pixels_row_30_24 = {data_out_rows[1105*col_length-1 -: col_length]};
assign pixels_col_30_25 = {data_out_cols[1106*col_length-1 -: col_length]};
assign pixels_row_30_25 = {data_out_rows[1106*col_length-1 -: col_length]};
assign pixels_col_30_26 = {data_out_cols[1107*col_length-1 -: col_length]};
assign pixels_row_30_26 = {data_out_rows[1107*col_length-1 -: col_length]};
assign pixels_col_30_27 = {data_out_cols[1108*col_length-1 -: col_length]};
assign pixels_row_30_27 = {data_out_rows[1108*col_length-1 -: col_length]};
assign pixels_col_30_28 = {data_out_cols[1109*col_length-1 -: col_length]};
assign pixels_row_30_28 = {data_out_rows[1109*col_length-1 -: col_length]};
assign pixels_col_30_29 = {data_out_cols[1110*col_length-1 -: col_length]};
assign pixels_row_30_29 = {data_out_rows[1110*col_length-1 -: col_length]};
assign pixels_col_30_30 = {data_out_cols[1111*col_length-1 -: col_length]};
assign pixels_row_30_30 = {data_out_rows[1111*col_length-1 -: col_length]};
assign pixels_col_30_31 = {data_out_cols[1112*col_length-1 -: col_length]};
assign pixels_row_30_31 = {data_out_rows[1112*col_length-1 -: col_length]};
assign pixels_col_30_32 = {data_out_cols[1113*col_length-1 -: col_length]};
assign pixels_row_30_32 = {data_out_rows[1113*col_length-1 -: col_length]};
assign pixels_col_30_33 = {data_out_cols[1114*col_length-1 -: col_length]};
assign pixels_row_30_33 = {data_out_rows[1114*col_length-1 -: col_length]};
assign pixels_col_30_34 = {data_out_cols[1115*col_length-1 -: col_length]};
assign pixels_row_30_34 = {data_out_rows[1115*col_length-1 -: col_length]};
assign pixels_col_30_35 = {data_out_cols[1116*col_length-1 -: col_length]};
assign pixels_row_30_35 = {data_out_rows[1116*col_length-1 -: col_length]};
assign pixels_col_31_0 = {data_out_cols[1117*col_length-1 -: col_length]};
assign pixels_row_31_0 = {data_out_rows[1117*col_length-1 -: col_length]};
assign pixels_col_31_1 = {data_out_cols[1118*col_length-1 -: col_length]};
assign pixels_row_31_1 = {data_out_rows[1118*col_length-1 -: col_length]};
assign pixels_col_31_2 = {data_out_cols[1119*col_length-1 -: col_length]};
assign pixels_row_31_2 = {data_out_rows[1119*col_length-1 -: col_length]};
assign pixels_col_31_3 = {data_out_cols[1120*col_length-1 -: col_length]};
assign pixels_row_31_3 = {data_out_rows[1120*col_length-1 -: col_length]};
assign pixels_col_31_4 = {data_out_cols[1121*col_length-1 -: col_length]};
assign pixels_row_31_4 = {data_out_rows[1121*col_length-1 -: col_length]};
assign pixels_col_31_5 = {data_out_cols[1122*col_length-1 -: col_length]};
assign pixels_row_31_5 = {data_out_rows[1122*col_length-1 -: col_length]};
assign pixels_col_31_6 = {data_out_cols[1123*col_length-1 -: col_length]};
assign pixels_row_31_6 = {data_out_rows[1123*col_length-1 -: col_length]};
assign pixels_col_31_7 = {data_out_cols[1124*col_length-1 -: col_length]};
assign pixels_row_31_7 = {data_out_rows[1124*col_length-1 -: col_length]};
assign pixels_col_31_8 = {data_out_cols[1125*col_length-1 -: col_length]};
assign pixels_row_31_8 = {data_out_rows[1125*col_length-1 -: col_length]};
assign pixels_col_31_9 = {data_out_cols[1126*col_length-1 -: col_length]};
assign pixels_row_31_9 = {data_out_rows[1126*col_length-1 -: col_length]};
assign pixels_col_31_10 = {data_out_cols[1127*col_length-1 -: col_length]};
assign pixels_row_31_10 = {data_out_rows[1127*col_length-1 -: col_length]};
assign pixels_col_31_11 = {data_out_cols[1128*col_length-1 -: col_length]};
assign pixels_row_31_11 = {data_out_rows[1128*col_length-1 -: col_length]};
assign pixels_col_31_12 = {data_out_cols[1129*col_length-1 -: col_length]};
assign pixels_row_31_12 = {data_out_rows[1129*col_length-1 -: col_length]};
assign pixels_col_31_13 = {data_out_cols[1130*col_length-1 -: col_length]};
assign pixels_row_31_13 = {data_out_rows[1130*col_length-1 -: col_length]};
assign pixels_col_31_14 = {data_out_cols[1131*col_length-1 -: col_length]};
assign pixels_row_31_14 = {data_out_rows[1131*col_length-1 -: col_length]};
assign pixels_col_31_15 = {data_out_cols[1132*col_length-1 -: col_length]};
assign pixels_row_31_15 = {data_out_rows[1132*col_length-1 -: col_length]};
assign pixels_col_31_16 = {data_out_cols[1133*col_length-1 -: col_length]};
assign pixels_row_31_16 = {data_out_rows[1133*col_length-1 -: col_length]};
assign pixels_col_31_17 = {data_out_cols[1134*col_length-1 -: col_length]};
assign pixels_row_31_17 = {data_out_rows[1134*col_length-1 -: col_length]};
assign pixels_col_31_18 = {data_out_cols[1135*col_length-1 -: col_length]};
assign pixels_row_31_18 = {data_out_rows[1135*col_length-1 -: col_length]};
assign pixels_col_31_19 = {data_out_cols[1136*col_length-1 -: col_length]};
assign pixels_row_31_19 = {data_out_rows[1136*col_length-1 -: col_length]};
assign pixels_col_31_20 = {data_out_cols[1137*col_length-1 -: col_length]};
assign pixels_row_31_20 = {data_out_rows[1137*col_length-1 -: col_length]};
assign pixels_col_31_21 = {data_out_cols[1138*col_length-1 -: col_length]};
assign pixels_row_31_21 = {data_out_rows[1138*col_length-1 -: col_length]};
assign pixels_col_31_22 = {data_out_cols[1139*col_length-1 -: col_length]};
assign pixels_row_31_22 = {data_out_rows[1139*col_length-1 -: col_length]};
assign pixels_col_31_23 = {data_out_cols[1140*col_length-1 -: col_length]};
assign pixels_row_31_23 = {data_out_rows[1140*col_length-1 -: col_length]};
assign pixels_col_31_24 = {data_out_cols[1141*col_length-1 -: col_length]};
assign pixels_row_31_24 = {data_out_rows[1141*col_length-1 -: col_length]};
assign pixels_col_31_25 = {data_out_cols[1142*col_length-1 -: col_length]};
assign pixels_row_31_25 = {data_out_rows[1142*col_length-1 -: col_length]};
assign pixels_col_31_26 = {data_out_cols[1143*col_length-1 -: col_length]};
assign pixels_row_31_26 = {data_out_rows[1143*col_length-1 -: col_length]};
assign pixels_col_31_27 = {data_out_cols[1144*col_length-1 -: col_length]};
assign pixels_row_31_27 = {data_out_rows[1144*col_length-1 -: col_length]};
assign pixels_col_31_28 = {data_out_cols[1145*col_length-1 -: col_length]};
assign pixels_row_31_28 = {data_out_rows[1145*col_length-1 -: col_length]};
assign pixels_col_31_29 = {data_out_cols[1146*col_length-1 -: col_length]};
assign pixels_row_31_29 = {data_out_rows[1146*col_length-1 -: col_length]};
assign pixels_col_31_30 = {data_out_cols[1147*col_length-1 -: col_length]};
assign pixels_row_31_30 = {data_out_rows[1147*col_length-1 -: col_length]};
assign pixels_col_31_31 = {data_out_cols[1148*col_length-1 -: col_length]};
assign pixels_row_31_31 = {data_out_rows[1148*col_length-1 -: col_length]};
assign pixels_col_31_32 = {data_out_cols[1149*col_length-1 -: col_length]};
assign pixels_row_31_32 = {data_out_rows[1149*col_length-1 -: col_length]};
assign pixels_col_31_33 = {data_out_cols[1150*col_length-1 -: col_length]};
assign pixels_row_31_33 = {data_out_rows[1150*col_length-1 -: col_length]};
assign pixels_col_31_34 = {data_out_cols[1151*col_length-1 -: col_length]};
assign pixels_row_31_34 = {data_out_rows[1151*col_length-1 -: col_length]};
assign pixels_col_31_35 = {data_out_cols[1152*col_length-1 -: col_length]};
assign pixels_row_31_35 = {data_out_rows[1152*col_length-1 -: col_length]};
assign pixels_col_32_0 = {data_out_cols[1153*col_length-1 -: col_length]};
assign pixels_row_32_0 = {data_out_rows[1153*col_length-1 -: col_length]};
assign pixels_col_32_1 = {data_out_cols[1154*col_length-1 -: col_length]};
assign pixels_row_32_1 = {data_out_rows[1154*col_length-1 -: col_length]};
assign pixels_col_32_2 = {data_out_cols[1155*col_length-1 -: col_length]};
assign pixels_row_32_2 = {data_out_rows[1155*col_length-1 -: col_length]};
assign pixels_col_32_3 = {data_out_cols[1156*col_length-1 -: col_length]};
assign pixels_row_32_3 = {data_out_rows[1156*col_length-1 -: col_length]};
assign pixels_col_32_4 = {data_out_cols[1157*col_length-1 -: col_length]};
assign pixels_row_32_4 = {data_out_rows[1157*col_length-1 -: col_length]};
assign pixels_col_32_5 = {data_out_cols[1158*col_length-1 -: col_length]};
assign pixels_row_32_5 = {data_out_rows[1158*col_length-1 -: col_length]};
assign pixels_col_32_6 = {data_out_cols[1159*col_length-1 -: col_length]};
assign pixels_row_32_6 = {data_out_rows[1159*col_length-1 -: col_length]};
assign pixels_col_32_7 = {data_out_cols[1160*col_length-1 -: col_length]};
assign pixels_row_32_7 = {data_out_rows[1160*col_length-1 -: col_length]};
assign pixels_col_32_8 = {data_out_cols[1161*col_length-1 -: col_length]};
assign pixels_row_32_8 = {data_out_rows[1161*col_length-1 -: col_length]};
assign pixels_col_32_9 = {data_out_cols[1162*col_length-1 -: col_length]};
assign pixels_row_32_9 = {data_out_rows[1162*col_length-1 -: col_length]};
assign pixels_col_32_10 = {data_out_cols[1163*col_length-1 -: col_length]};
assign pixels_row_32_10 = {data_out_rows[1163*col_length-1 -: col_length]};
assign pixels_col_32_11 = {data_out_cols[1164*col_length-1 -: col_length]};
assign pixels_row_32_11 = {data_out_rows[1164*col_length-1 -: col_length]};
assign pixels_col_32_12 = {data_out_cols[1165*col_length-1 -: col_length]};
assign pixels_row_32_12 = {data_out_rows[1165*col_length-1 -: col_length]};
assign pixels_col_32_13 = {data_out_cols[1166*col_length-1 -: col_length]};
assign pixels_row_32_13 = {data_out_rows[1166*col_length-1 -: col_length]};
assign pixels_col_32_14 = {data_out_cols[1167*col_length-1 -: col_length]};
assign pixels_row_32_14 = {data_out_rows[1167*col_length-1 -: col_length]};
assign pixels_col_32_15 = {data_out_cols[1168*col_length-1 -: col_length]};
assign pixels_row_32_15 = {data_out_rows[1168*col_length-1 -: col_length]};
assign pixels_col_32_16 = {data_out_cols[1169*col_length-1 -: col_length]};
assign pixels_row_32_16 = {data_out_rows[1169*col_length-1 -: col_length]};
assign pixels_col_32_17 = {data_out_cols[1170*col_length-1 -: col_length]};
assign pixels_row_32_17 = {data_out_rows[1170*col_length-1 -: col_length]};
assign pixels_col_32_18 = {data_out_cols[1171*col_length-1 -: col_length]};
assign pixels_row_32_18 = {data_out_rows[1171*col_length-1 -: col_length]};
assign pixels_col_32_19 = {data_out_cols[1172*col_length-1 -: col_length]};
assign pixels_row_32_19 = {data_out_rows[1172*col_length-1 -: col_length]};
assign pixels_col_32_20 = {data_out_cols[1173*col_length-1 -: col_length]};
assign pixels_row_32_20 = {data_out_rows[1173*col_length-1 -: col_length]};
assign pixels_col_32_21 = {data_out_cols[1174*col_length-1 -: col_length]};
assign pixels_row_32_21 = {data_out_rows[1174*col_length-1 -: col_length]};
assign pixels_col_32_22 = {data_out_cols[1175*col_length-1 -: col_length]};
assign pixels_row_32_22 = {data_out_rows[1175*col_length-1 -: col_length]};
assign pixels_col_32_23 = {data_out_cols[1176*col_length-1 -: col_length]};
assign pixels_row_32_23 = {data_out_rows[1176*col_length-1 -: col_length]};
assign pixels_col_32_24 = {data_out_cols[1177*col_length-1 -: col_length]};
assign pixels_row_32_24 = {data_out_rows[1177*col_length-1 -: col_length]};
assign pixels_col_32_25 = {data_out_cols[1178*col_length-1 -: col_length]};
assign pixels_row_32_25 = {data_out_rows[1178*col_length-1 -: col_length]};
assign pixels_col_32_26 = {data_out_cols[1179*col_length-1 -: col_length]};
assign pixels_row_32_26 = {data_out_rows[1179*col_length-1 -: col_length]};
assign pixels_col_32_27 = {data_out_cols[1180*col_length-1 -: col_length]};
assign pixels_row_32_27 = {data_out_rows[1180*col_length-1 -: col_length]};
assign pixels_col_32_28 = {data_out_cols[1181*col_length-1 -: col_length]};
assign pixels_row_32_28 = {data_out_rows[1181*col_length-1 -: col_length]};
assign pixels_col_32_29 = {data_out_cols[1182*col_length-1 -: col_length]};
assign pixels_row_32_29 = {data_out_rows[1182*col_length-1 -: col_length]};
assign pixels_col_32_30 = {data_out_cols[1183*col_length-1 -: col_length]};
assign pixels_row_32_30 = {data_out_rows[1183*col_length-1 -: col_length]};
assign pixels_col_32_31 = {data_out_cols[1184*col_length-1 -: col_length]};
assign pixels_row_32_31 = {data_out_rows[1184*col_length-1 -: col_length]};
assign pixels_col_32_32 = {data_out_cols[1185*col_length-1 -: col_length]};
assign pixels_row_32_32 = {data_out_rows[1185*col_length-1 -: col_length]};
assign pixels_col_32_33 = {data_out_cols[1186*col_length-1 -: col_length]};
assign pixels_row_32_33 = {data_out_rows[1186*col_length-1 -: col_length]};
assign pixels_col_32_34 = {data_out_cols[1187*col_length-1 -: col_length]};
assign pixels_row_32_34 = {data_out_rows[1187*col_length-1 -: col_length]};
assign pixels_col_32_35 = {data_out_cols[1188*col_length-1 -: col_length]};
assign pixels_row_32_35 = {data_out_rows[1188*col_length-1 -: col_length]};
assign pixels_col_33_0 = {data_out_cols[1189*col_length-1 -: col_length]};
assign pixels_row_33_0 = {data_out_rows[1189*col_length-1 -: col_length]};
assign pixels_col_33_1 = {data_out_cols[1190*col_length-1 -: col_length]};
assign pixels_row_33_1 = {data_out_rows[1190*col_length-1 -: col_length]};
assign pixels_col_33_2 = {data_out_cols[1191*col_length-1 -: col_length]};
assign pixels_row_33_2 = {data_out_rows[1191*col_length-1 -: col_length]};
assign pixels_col_33_3 = {data_out_cols[1192*col_length-1 -: col_length]};
assign pixels_row_33_3 = {data_out_rows[1192*col_length-1 -: col_length]};
assign pixels_col_33_4 = {data_out_cols[1193*col_length-1 -: col_length]};
assign pixels_row_33_4 = {data_out_rows[1193*col_length-1 -: col_length]};
assign pixels_col_33_5 = {data_out_cols[1194*col_length-1 -: col_length]};
assign pixels_row_33_5 = {data_out_rows[1194*col_length-1 -: col_length]};
assign pixels_col_33_6 = {data_out_cols[1195*col_length-1 -: col_length]};
assign pixels_row_33_6 = {data_out_rows[1195*col_length-1 -: col_length]};
assign pixels_col_33_7 = {data_out_cols[1196*col_length-1 -: col_length]};
assign pixels_row_33_7 = {data_out_rows[1196*col_length-1 -: col_length]};
assign pixels_col_33_8 = {data_out_cols[1197*col_length-1 -: col_length]};
assign pixels_row_33_8 = {data_out_rows[1197*col_length-1 -: col_length]};
assign pixels_col_33_9 = {data_out_cols[1198*col_length-1 -: col_length]};
assign pixels_row_33_9 = {data_out_rows[1198*col_length-1 -: col_length]};
assign pixels_col_33_10 = {data_out_cols[1199*col_length-1 -: col_length]};
assign pixels_row_33_10 = {data_out_rows[1199*col_length-1 -: col_length]};
assign pixels_col_33_11 = {data_out_cols[1200*col_length-1 -: col_length]};
assign pixels_row_33_11 = {data_out_rows[1200*col_length-1 -: col_length]};
assign pixels_col_33_12 = {data_out_cols[1201*col_length-1 -: col_length]};
assign pixels_row_33_12 = {data_out_rows[1201*col_length-1 -: col_length]};
assign pixels_col_33_13 = {data_out_cols[1202*col_length-1 -: col_length]};
assign pixels_row_33_13 = {data_out_rows[1202*col_length-1 -: col_length]};
assign pixels_col_33_14 = {data_out_cols[1203*col_length-1 -: col_length]};
assign pixels_row_33_14 = {data_out_rows[1203*col_length-1 -: col_length]};
assign pixels_col_33_15 = {data_out_cols[1204*col_length-1 -: col_length]};
assign pixels_row_33_15 = {data_out_rows[1204*col_length-1 -: col_length]};
assign pixels_col_33_16 = {data_out_cols[1205*col_length-1 -: col_length]};
assign pixels_row_33_16 = {data_out_rows[1205*col_length-1 -: col_length]};
assign pixels_col_33_17 = {data_out_cols[1206*col_length-1 -: col_length]};
assign pixels_row_33_17 = {data_out_rows[1206*col_length-1 -: col_length]};
assign pixels_col_33_18 = {data_out_cols[1207*col_length-1 -: col_length]};
assign pixels_row_33_18 = {data_out_rows[1207*col_length-1 -: col_length]};
assign pixels_col_33_19 = {data_out_cols[1208*col_length-1 -: col_length]};
assign pixels_row_33_19 = {data_out_rows[1208*col_length-1 -: col_length]};
assign pixels_col_33_20 = {data_out_cols[1209*col_length-1 -: col_length]};
assign pixels_row_33_20 = {data_out_rows[1209*col_length-1 -: col_length]};
assign pixels_col_33_21 = {data_out_cols[1210*col_length-1 -: col_length]};
assign pixels_row_33_21 = {data_out_rows[1210*col_length-1 -: col_length]};
assign pixels_col_33_22 = {data_out_cols[1211*col_length-1 -: col_length]};
assign pixels_row_33_22 = {data_out_rows[1211*col_length-1 -: col_length]};
assign pixels_col_33_23 = {data_out_cols[1212*col_length-1 -: col_length]};
assign pixels_row_33_23 = {data_out_rows[1212*col_length-1 -: col_length]};
assign pixels_col_33_24 = {data_out_cols[1213*col_length-1 -: col_length]};
assign pixels_row_33_24 = {data_out_rows[1213*col_length-1 -: col_length]};
assign pixels_col_33_25 = {data_out_cols[1214*col_length-1 -: col_length]};
assign pixels_row_33_25 = {data_out_rows[1214*col_length-1 -: col_length]};
assign pixels_col_33_26 = {data_out_cols[1215*col_length-1 -: col_length]};
assign pixels_row_33_26 = {data_out_rows[1215*col_length-1 -: col_length]};
assign pixels_col_33_27 = {data_out_cols[1216*col_length-1 -: col_length]};
assign pixels_row_33_27 = {data_out_rows[1216*col_length-1 -: col_length]};
assign pixels_col_33_28 = {data_out_cols[1217*col_length-1 -: col_length]};
assign pixels_row_33_28 = {data_out_rows[1217*col_length-1 -: col_length]};
assign pixels_col_33_29 = {data_out_cols[1218*col_length-1 -: col_length]};
assign pixels_row_33_29 = {data_out_rows[1218*col_length-1 -: col_length]};
assign pixels_col_33_30 = {data_out_cols[1219*col_length-1 -: col_length]};
assign pixels_row_33_30 = {data_out_rows[1219*col_length-1 -: col_length]};
assign pixels_col_33_31 = {data_out_cols[1220*col_length-1 -: col_length]};
assign pixels_row_33_31 = {data_out_rows[1220*col_length-1 -: col_length]};
assign pixels_col_33_32 = {data_out_cols[1221*col_length-1 -: col_length]};
assign pixels_row_33_32 = {data_out_rows[1221*col_length-1 -: col_length]};
assign pixels_col_33_33 = {data_out_cols[1222*col_length-1 -: col_length]};
assign pixels_row_33_33 = {data_out_rows[1222*col_length-1 -: col_length]};
assign pixels_col_33_34 = {data_out_cols[1223*col_length-1 -: col_length]};
assign pixels_row_33_34 = {data_out_rows[1223*col_length-1 -: col_length]};
assign pixels_col_33_35 = {data_out_cols[1224*col_length-1 -: col_length]};
assign pixels_row_33_35 = {data_out_rows[1224*col_length-1 -: col_length]};
assign pixels_col_34_0 = {data_out_cols[1225*col_length-1 -: col_length]};
assign pixels_row_34_0 = {data_out_rows[1225*col_length-1 -: col_length]};
assign pixels_col_34_1 = {data_out_cols[1226*col_length-1 -: col_length]};
assign pixels_row_34_1 = {data_out_rows[1226*col_length-1 -: col_length]};
assign pixels_col_34_2 = {data_out_cols[1227*col_length-1 -: col_length]};
assign pixels_row_34_2 = {data_out_rows[1227*col_length-1 -: col_length]};
assign pixels_col_34_3 = {data_out_cols[1228*col_length-1 -: col_length]};
assign pixels_row_34_3 = {data_out_rows[1228*col_length-1 -: col_length]};
assign pixels_col_34_4 = {data_out_cols[1229*col_length-1 -: col_length]};
assign pixels_row_34_4 = {data_out_rows[1229*col_length-1 -: col_length]};
assign pixels_col_34_5 = {data_out_cols[1230*col_length-1 -: col_length]};
assign pixels_row_34_5 = {data_out_rows[1230*col_length-1 -: col_length]};
assign pixels_col_34_6 = {data_out_cols[1231*col_length-1 -: col_length]};
assign pixels_row_34_6 = {data_out_rows[1231*col_length-1 -: col_length]};
assign pixels_col_34_7 = {data_out_cols[1232*col_length-1 -: col_length]};
assign pixels_row_34_7 = {data_out_rows[1232*col_length-1 -: col_length]};
assign pixels_col_34_8 = {data_out_cols[1233*col_length-1 -: col_length]};
assign pixels_row_34_8 = {data_out_rows[1233*col_length-1 -: col_length]};
assign pixels_col_34_9 = {data_out_cols[1234*col_length-1 -: col_length]};
assign pixels_row_34_9 = {data_out_rows[1234*col_length-1 -: col_length]};
assign pixels_col_34_10 = {data_out_cols[1235*col_length-1 -: col_length]};
assign pixels_row_34_10 = {data_out_rows[1235*col_length-1 -: col_length]};
assign pixels_col_34_11 = {data_out_cols[1236*col_length-1 -: col_length]};
assign pixels_row_34_11 = {data_out_rows[1236*col_length-1 -: col_length]};
assign pixels_col_34_12 = {data_out_cols[1237*col_length-1 -: col_length]};
assign pixels_row_34_12 = {data_out_rows[1237*col_length-1 -: col_length]};
assign pixels_col_34_13 = {data_out_cols[1238*col_length-1 -: col_length]};
assign pixels_row_34_13 = {data_out_rows[1238*col_length-1 -: col_length]};
assign pixels_col_34_14 = {data_out_cols[1239*col_length-1 -: col_length]};
assign pixels_row_34_14 = {data_out_rows[1239*col_length-1 -: col_length]};
assign pixels_col_34_15 = {data_out_cols[1240*col_length-1 -: col_length]};
assign pixels_row_34_15 = {data_out_rows[1240*col_length-1 -: col_length]};
assign pixels_col_34_16 = {data_out_cols[1241*col_length-1 -: col_length]};
assign pixels_row_34_16 = {data_out_rows[1241*col_length-1 -: col_length]};
assign pixels_col_34_17 = {data_out_cols[1242*col_length-1 -: col_length]};
assign pixels_row_34_17 = {data_out_rows[1242*col_length-1 -: col_length]};
assign pixels_col_34_18 = {data_out_cols[1243*col_length-1 -: col_length]};
assign pixels_row_34_18 = {data_out_rows[1243*col_length-1 -: col_length]};
assign pixels_col_34_19 = {data_out_cols[1244*col_length-1 -: col_length]};
assign pixels_row_34_19 = {data_out_rows[1244*col_length-1 -: col_length]};
assign pixels_col_34_20 = {data_out_cols[1245*col_length-1 -: col_length]};
assign pixels_row_34_20 = {data_out_rows[1245*col_length-1 -: col_length]};
assign pixels_col_34_21 = {data_out_cols[1246*col_length-1 -: col_length]};
assign pixels_row_34_21 = {data_out_rows[1246*col_length-1 -: col_length]};
assign pixels_col_34_22 = {data_out_cols[1247*col_length-1 -: col_length]};
assign pixels_row_34_22 = {data_out_rows[1247*col_length-1 -: col_length]};
assign pixels_col_34_23 = {data_out_cols[1248*col_length-1 -: col_length]};
assign pixels_row_34_23 = {data_out_rows[1248*col_length-1 -: col_length]};
assign pixels_col_34_24 = {data_out_cols[1249*col_length-1 -: col_length]};
assign pixels_row_34_24 = {data_out_rows[1249*col_length-1 -: col_length]};
assign pixels_col_34_25 = {data_out_cols[1250*col_length-1 -: col_length]};
assign pixels_row_34_25 = {data_out_rows[1250*col_length-1 -: col_length]};
assign pixels_col_34_26 = {data_out_cols[1251*col_length-1 -: col_length]};
assign pixels_row_34_26 = {data_out_rows[1251*col_length-1 -: col_length]};
assign pixels_col_34_27 = {data_out_cols[1252*col_length-1 -: col_length]};
assign pixels_row_34_27 = {data_out_rows[1252*col_length-1 -: col_length]};
assign pixels_col_34_28 = {data_out_cols[1253*col_length-1 -: col_length]};
assign pixels_row_34_28 = {data_out_rows[1253*col_length-1 -: col_length]};
assign pixels_col_34_29 = {data_out_cols[1254*col_length-1 -: col_length]};
assign pixels_row_34_29 = {data_out_rows[1254*col_length-1 -: col_length]};
assign pixels_col_34_30 = {data_out_cols[1255*col_length-1 -: col_length]};
assign pixels_row_34_30 = {data_out_rows[1255*col_length-1 -: col_length]};
assign pixels_col_34_31 = {data_out_cols[1256*col_length-1 -: col_length]};
assign pixels_row_34_31 = {data_out_rows[1256*col_length-1 -: col_length]};
assign pixels_col_34_32 = {data_out_cols[1257*col_length-1 -: col_length]};
assign pixels_row_34_32 = {data_out_rows[1257*col_length-1 -: col_length]};
assign pixels_col_34_33 = {data_out_cols[1258*col_length-1 -: col_length]};
assign pixels_row_34_33 = {data_out_rows[1258*col_length-1 -: col_length]};
assign pixels_col_34_34 = {data_out_cols[1259*col_length-1 -: col_length]};
assign pixels_row_34_34 = {data_out_rows[1259*col_length-1 -: col_length]};
assign pixels_col_34_35 = {data_out_cols[1260*col_length-1 -: col_length]};
assign pixels_row_34_35 = {data_out_rows[1260*col_length-1 -: col_length]};
assign pixels_col_35_0 = {data_out_cols[1261*col_length-1 -: col_length]};
assign pixels_row_35_0 = {data_out_rows[1261*col_length-1 -: col_length]};
assign pixels_col_35_1 = {data_out_cols[1262*col_length-1 -: col_length]};
assign pixels_row_35_1 = {data_out_rows[1262*col_length-1 -: col_length]};
assign pixels_col_35_2 = {data_out_cols[1263*col_length-1 -: col_length]};
assign pixels_row_35_2 = {data_out_rows[1263*col_length-1 -: col_length]};
assign pixels_col_35_3 = {data_out_cols[1264*col_length-1 -: col_length]};
assign pixels_row_35_3 = {data_out_rows[1264*col_length-1 -: col_length]};
assign pixels_col_35_4 = {data_out_cols[1265*col_length-1 -: col_length]};
assign pixels_row_35_4 = {data_out_rows[1265*col_length-1 -: col_length]};
assign pixels_col_35_5 = {data_out_cols[1266*col_length-1 -: col_length]};
assign pixels_row_35_5 = {data_out_rows[1266*col_length-1 -: col_length]};
assign pixels_col_35_6 = {data_out_cols[1267*col_length-1 -: col_length]};
assign pixels_row_35_6 = {data_out_rows[1267*col_length-1 -: col_length]};
assign pixels_col_35_7 = {data_out_cols[1268*col_length-1 -: col_length]};
assign pixels_row_35_7 = {data_out_rows[1268*col_length-1 -: col_length]};
assign pixels_col_35_8 = {data_out_cols[1269*col_length-1 -: col_length]};
assign pixels_row_35_8 = {data_out_rows[1269*col_length-1 -: col_length]};
assign pixels_col_35_9 = {data_out_cols[1270*col_length-1 -: col_length]};
assign pixels_row_35_9 = {data_out_rows[1270*col_length-1 -: col_length]};
assign pixels_col_35_10 = {data_out_cols[1271*col_length-1 -: col_length]};
assign pixels_row_35_10 = {data_out_rows[1271*col_length-1 -: col_length]};
assign pixels_col_35_11 = {data_out_cols[1272*col_length-1 -: col_length]};
assign pixels_row_35_11 = {data_out_rows[1272*col_length-1 -: col_length]};
assign pixels_col_35_12 = {data_out_cols[1273*col_length-1 -: col_length]};
assign pixels_row_35_12 = {data_out_rows[1273*col_length-1 -: col_length]};
assign pixels_col_35_13 = {data_out_cols[1274*col_length-1 -: col_length]};
assign pixels_row_35_13 = {data_out_rows[1274*col_length-1 -: col_length]};
assign pixels_col_35_14 = {data_out_cols[1275*col_length-1 -: col_length]};
assign pixels_row_35_14 = {data_out_rows[1275*col_length-1 -: col_length]};
assign pixels_col_35_15 = {data_out_cols[1276*col_length-1 -: col_length]};
assign pixels_row_35_15 = {data_out_rows[1276*col_length-1 -: col_length]};
assign pixels_col_35_16 = {data_out_cols[1277*col_length-1 -: col_length]};
assign pixels_row_35_16 = {data_out_rows[1277*col_length-1 -: col_length]};
assign pixels_col_35_17 = {data_out_cols[1278*col_length-1 -: col_length]};
assign pixels_row_35_17 = {data_out_rows[1278*col_length-1 -: col_length]};
assign pixels_col_35_18 = {data_out_cols[1279*col_length-1 -: col_length]};
assign pixels_row_35_18 = {data_out_rows[1279*col_length-1 -: col_length]};
assign pixels_col_35_19 = {data_out_cols[1280*col_length-1 -: col_length]};
assign pixels_row_35_19 = {data_out_rows[1280*col_length-1 -: col_length]};
assign pixels_col_35_20 = {data_out_cols[1281*col_length-1 -: col_length]};
assign pixels_row_35_20 = {data_out_rows[1281*col_length-1 -: col_length]};
assign pixels_col_35_21 = {data_out_cols[1282*col_length-1 -: col_length]};
assign pixels_row_35_21 = {data_out_rows[1282*col_length-1 -: col_length]};
assign pixels_col_35_22 = {data_out_cols[1283*col_length-1 -: col_length]};
assign pixels_row_35_22 = {data_out_rows[1283*col_length-1 -: col_length]};
assign pixels_col_35_23 = {data_out_cols[1284*col_length-1 -: col_length]};
assign pixels_row_35_23 = {data_out_rows[1284*col_length-1 -: col_length]};
assign pixels_col_35_24 = {data_out_cols[1285*col_length-1 -: col_length]};
assign pixels_row_35_24 = {data_out_rows[1285*col_length-1 -: col_length]};
assign pixels_col_35_25 = {data_out_cols[1286*col_length-1 -: col_length]};
assign pixels_row_35_25 = {data_out_rows[1286*col_length-1 -: col_length]};
assign pixels_col_35_26 = {data_out_cols[1287*col_length-1 -: col_length]};
assign pixels_row_35_26 = {data_out_rows[1287*col_length-1 -: col_length]};
assign pixels_col_35_27 = {data_out_cols[1288*col_length-1 -: col_length]};
assign pixels_row_35_27 = {data_out_rows[1288*col_length-1 -: col_length]};
assign pixels_col_35_28 = {data_out_cols[1289*col_length-1 -: col_length]};
assign pixels_row_35_28 = {data_out_rows[1289*col_length-1 -: col_length]};
assign pixels_col_35_29 = {data_out_cols[1290*col_length-1 -: col_length]};
assign pixels_row_35_29 = {data_out_rows[1290*col_length-1 -: col_length]};
assign pixels_col_35_30 = {data_out_cols[1291*col_length-1 -: col_length]};
assign pixels_row_35_30 = {data_out_rows[1291*col_length-1 -: col_length]};
assign pixels_col_35_31 = {data_out_cols[1292*col_length-1 -: col_length]};
assign pixels_row_35_31 = {data_out_rows[1292*col_length-1 -: col_length]};
assign pixels_col_35_32 = {data_out_cols[1293*col_length-1 -: col_length]};
assign pixels_row_35_32 = {data_out_rows[1293*col_length-1 -: col_length]};
assign pixels_col_35_33 = {data_out_cols[1294*col_length-1 -: col_length]};
assign pixels_row_35_33 = {data_out_rows[1294*col_length-1 -: col_length]};
assign pixels_col_35_34 = {data_out_cols[1295*col_length-1 -: col_length]};
assign pixels_row_35_34 = {data_out_rows[1295*col_length-1 -: col_length]};
assign pixels_col_35_35 = {data_out_cols[1296*col_length-1 -: col_length]};
assign pixels_row_35_35 = {data_out_rows[1296*col_length-1 -: col_length]};
//iter
integer i;

initial begin
    #0      rst = 0;
            clk = 1;
    #10     rst = 1;
            data_in = 0;
    #10     rst = 0;
    #100    in_valid = 1;
            for (i=0;i<(image_size*image_size);i=i+1)begin
                data_in[word_length-1:0] = {pe_input_feature_value[(i+1)*word_length-1 -:word_length]};
                //data_in[word_length-1:0] = i+1;
                #10;
            end
    #1000;
    

    $finish;
    
end




always #5 clk = ~clk;
CSR#
(
    .col_length(col_length), 
    .word_length(word_length), 
    .double_word_length(double_word_length), 
    .kernel_size(kernel_size), 
    .image_size(image_size)
)u1
(
    .clk(clk), 
    .rst(rst), 
    .in_valid(in_valid),
    .data_in(data_in),
    .data_out(data_out),
    .data_out_cols(data_out_cols),
    .data_out_rows(data_out_rows)
);



endmodule