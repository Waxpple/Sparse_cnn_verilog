`timescale 1ns/1ns
module conv_tb();
parameter col_length = 8;
parameter word_length = 8;
parameter double_word_length = 16;
parameter kernel_size = 5;
parameter image_size = 36;

reg clk;
reg rst;
reg signed [word_length-1:0] data_in;
reg in_valid;
reg [10368-1 :0] pe_input_feature_value='h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_f0_dd_39_f3_f7_06_02_f7_02_f6_fc_15_f9_ff_15_08_fe_fb_f0_01_e5_09_00_f9_1d_fa_f6_ec_00_00_00_00_00_00_00_00_fd_f2_fb_f2_eb_f3_fa_f3_12_fc_f8_0b_03_fe_f1_f6_07_f7_eb_0a_17_f5_05_01_18_1f_f1_09_00_00_00_00_00_00_00_00_07_04_f3_0c_fa_f6_01_0d_07_e5_06_f8_0e_0b_f9_03_fc_e1_0b_f2_15_fa_0d_ee_08_f9_ed_ff_00_00_00_00_00_00_00_00_f8_fc_fa_f8_e8_07_f2_0f_00_da_08_fb_03_06_f2_f0_07_03_06_fb_e9_f5_13_06_fa_0d_05_0a_00_00_00_00_00_00_00_00_f1_0d_f6_03_fa_03_17_1c_06_e4_13_03_11_0c_f4_15_fb_0d_fd_07_02_0b_f5_0e_ea_e0_ee_04_00_00_00_00_00_00_00_00_f2_fb_01_01_e7_01_ea_07_0e_fc_08_1f_1a_04_fa_ef_02_00_d8_fa_eb_ee_0d_f1_f4_ff_01_fd_00_00_00_00_00_00_00_00_18_eb_f2_08_12_04_0b_fb_f7_0a_00_0b_05_f7_f2_0a_1a_e6_15_0e_29_12_f8_08_dd_f9_0f_10_00_00_00_00_00_00_00_00_05_df_02_07_f1_fe_01_0c_dc_fb_fb_fb_16_15_e8_f8_02_fe_0e_10_0d_fb_fa_02_fd_e5_03_09_00_00_00_00_00_00_00_00_f5_f9_fd_e5_05_0a_03_04_0c_0a_1d_0f_0e_1b_fb_26_f2_ec_08_08_f8_03_08_1b_fc_19_f7_f4_00_00_00_00_00_00_00_00_13_00_fc_13_00_1e_12_fc_11_15_11_00_f7_dd_f6_05_0d_f3_1a_13_fd_18_0e_f1_14_09_dd_0a_00_00_00_00_00_00_00_00_ed_e6_f1_06_ed_fc_fb_fe_10_07_f0_17_15_03_07_f5_0a_13_06_13_fa_1c_07_05_03_ee_eb_f1_00_00_00_00_00_00_00_00_dc_09_f6_fc_fb_04_d9_f9_08_01_08_18_15_25_e6_fe_f9_03_f1_fc_f3_fb_0e_00_f2_f0_0a_f7_00_00_00_00_00_00_00_00_06_0b_f8_26_f5_0c_e6_09_f7_fe_fa_04_fa_0b_dc_f8_12_e4_f3_f5_02_0a_f9_20_fd_04_12_fa_00_00_00_00_00_00_00_00_fb_03_15_e2_ef_f4_01_19_0c_fd_fc_fc_03_0f_18_f2_05_e9_f2_22_04_ef_f5_03_fd_10_f4_e2_00_00_00_00_00_00_00_00_0b_07_02_ec_f8_01_0e_fe_fc_03_ef_eb_f1_f9_04_06_09_15_fc_01_03_f9_0d_ec_f2_2a_e9_01_00_00_00_00_00_00_00_00_0b_12_e9_ff_e9_0d_f3_0f_e4_02_08_0d_e9_e3_fc_05_f3_f6_fd_ee_fc_e4_f5_f3_ef_e1_06_f5_00_00_00_00_00_00_00_00_0b_00_16_e1_f2_f1_06_03_ff_fa_07_f3_09_f7_0a_0a_0c_ff_1f_f4_0f_ef_fb_15_02_e6_fd_f9_00_00_00_00_00_00_00_00_08_f1_ff_f1_eb_11_f4_ea_fd_f3_f0_05_0a_e9_05_0a_f7_e8_f7_f2_11_f4_03_f5_13_e9_fb_fc_00_00_00_00_00_00_00_00_04_fb_0a_01_f9_04_00_03_f7_fb_0b_2c_13_0a_10_ec_08_eb_17_fa_1e_05_18_f4_02_01_0a_03_00_00_00_00_00_00_00_00_ff_02_f6_f9_f6_00_07_01_01_f2_0d_19_fc_05_ef_f3_0c_e7_0d_e1_07_09_26_ff_f8_0a_cf_f1_00_00_00_00_00_00_00_00_e9_08_04_ff_fe_e4_dc_fa_05_fc_23_09_ff_03_09_04_18_1a_f4_02_d7_2a_ed_09_07_14_f0_ff_00_00_00_00_00_00_00_00_0f_09_0f_f8_08_f1_21_02_27_fc_f8_fb_ef_11_ee_f9_17_13_01_2c_04_f6_1c_e8_f7_f8_fa_08_00_00_00_00_00_00_00_00_13_f6_11_24_fb_00_f4_09_0d_ff_ff_2c_f2_0f_2b_e0_fa_0c_04_25_fa_0a_0c_0c_15_f9_07_f6_00_00_00_00_00_00_00_00_fa_f7_07_20_f8_17_10_07_0a_07_1a_04_0b_f6_ff_1a_ef_e6_03_02_06_1f_fb_0c_06_f9_ff_04_00_00_00_00_00_00_00_00_1c_ec_f8_09_fc_20_e8_0e_f6_ed_f6_1c_00_e9_f6_07_15_f1_06_12_f9_e7_ef_08_ed_fb_16_fd_00_00_00_00_00_00_00_00_13_0d_fa_df_f0_09_e6_fd_f5_09_03_fa_17_fa_2f_16_ff_09_10_04_09_fe_fd_0d_f6_f2_e3_e2_00_00_00_00_00_00_00_00_f1_12_1b_ed_fb_18_fe_fd_01_1b_01_01_f3_1d_ff_07_0f_fe_05_ef_ef_38_fc_fb_ee_fc_f0_0e_00_00_00_00_00_00_00_00_02_37_0c_f4_1e_e1_04_f4_f4_0a_22_06_01_f0_00_00_1d_0d_fd_1f_f4_06_02_fe_07_ec_12_f7_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;

wire out_valid;
reg [kernel_size*kernel_size*word_length-1 :0] weight_value;
wire signed  [word_length*2-1:0] pixels_0_0, pixels_0_1, pixels_0_2, pixels_0_3, pixels_0_4, pixels_0_5, pixels_0_6, pixels_0_7, pixels_0_8, pixels_0_9, pixels_0_10, pixels_0_11, pixels_0_12, pixels_0_13, pixels_0_14, pixels_0_15, pixels_0_16, pixels_0_17, pixels_0_18, pixels_0_19, pixels_0_20, pixels_0_21, pixels_0_22, pixels_0_23, pixels_0_24, pixels_0_25, pixels_0_26, pixels_0_27, pixels_0_28, pixels_0_29, pixels_0_30, pixels_0_31, pixels_1_0, pixels_1_1, pixels_1_2, pixels_1_3, pixels_1_4, pixels_1_5, pixels_1_6, pixels_1_7, pixels_1_8, pixels_1_9, pixels_1_10, pixels_1_11, pixels_1_12, pixels_1_13, pixels_1_14, pixels_1_15, pixels_1_16, pixels_1_17, pixels_1_18, pixels_1_19, pixels_1_20, pixels_1_21, pixels_1_22, pixels_1_23, pixels_1_24, pixels_1_25, pixels_1_26, pixels_1_27, pixels_1_28, pixels_1_29, pixels_1_30, pixels_1_31, pixels_2_0, pixels_2_1, pixels_2_2, pixels_2_3, pixels_2_4, pixels_2_5, pixels_2_6, pixels_2_7, pixels_2_8, pixels_2_9, pixels_2_10, pixels_2_11, pixels_2_12, pixels_2_13, pixels_2_14, pixels_2_15, pixels_2_16, pixels_2_17, pixels_2_18, pixels_2_19, pixels_2_20, pixels_2_21, pixels_2_22, pixels_2_23, pixels_2_24, pixels_2_25, pixels_2_26, pixels_2_27, pixels_2_28, pixels_2_29, pixels_2_30, pixels_2_31, pixels_3_0, pixels_3_1, pixels_3_2, pixels_3_3, pixels_3_4, pixels_3_5, pixels_3_6, pixels_3_7, pixels_3_8, pixels_3_9, pixels_3_10, pixels_3_11, pixels_3_12, pixels_3_13, pixels_3_14, pixels_3_15, pixels_3_16, pixels_3_17, pixels_3_18, pixels_3_19, pixels_3_20, pixels_3_21, pixels_3_22, pixels_3_23, pixels_3_24, pixels_3_25, pixels_3_26, pixels_3_27, pixels_3_28, pixels_3_29, pixels_3_30, pixels_3_31, pixels_4_0, pixels_4_1, pixels_4_2, pixels_4_3, pixels_4_4, pixels_4_5, pixels_4_6, pixels_4_7, pixels_4_8, pixels_4_9, pixels_4_10, pixels_4_11, pixels_4_12, pixels_4_13, pixels_4_14, pixels_4_15, pixels_4_16, pixels_4_17, pixels_4_18, pixels_4_19, pixels_4_20, pixels_4_21, pixels_4_22, pixels_4_23, pixels_4_24, pixels_4_25, pixels_4_26, pixels_4_27, pixels_4_28, pixels_4_29, pixels_4_30, pixels_4_31, pixels_5_0, pixels_5_1, pixels_5_2, pixels_5_3, pixels_5_4, pixels_5_5, pixels_5_6, pixels_5_7, pixels_5_8, pixels_5_9, pixels_5_10, pixels_5_11, pixels_5_12, pixels_5_13, pixels_5_14, pixels_5_15, pixels_5_16, pixels_5_17, pixels_5_18, pixels_5_19, pixels_5_20, pixels_5_21, pixels_5_22, pixels_5_23, pixels_5_24, pixels_5_25, pixels_5_26, pixels_5_27, pixels_5_28, pixels_5_29, pixels_5_30, pixels_5_31, pixels_6_0, pixels_6_1, pixels_6_2, pixels_6_3, pixels_6_4, pixels_6_5, pixels_6_6, pixels_6_7, pixels_6_8, pixels_6_9, pixels_6_10, pixels_6_11, pixels_6_12, pixels_6_13, pixels_6_14, pixels_6_15, pixels_6_16, pixels_6_17, pixels_6_18, pixels_6_19, pixels_6_20, pixels_6_21, pixels_6_22, pixels_6_23, pixels_6_24, pixels_6_25, pixels_6_26, pixels_6_27, pixels_6_28, pixels_6_29, pixels_6_30, pixels_6_31, pixels_7_0, pixels_7_1, pixels_7_2, pixels_7_3, pixels_7_4, pixels_7_5, pixels_7_6, pixels_7_7, pixels_7_8, pixels_7_9, pixels_7_10, pixels_7_11, pixels_7_12, pixels_7_13, pixels_7_14, pixels_7_15, pixels_7_16, pixels_7_17, pixels_7_18, pixels_7_19, pixels_7_20, pixels_7_21, pixels_7_22, pixels_7_23, pixels_7_24, pixels_7_25, pixels_7_26, pixels_7_27, pixels_7_28, pixels_7_29, pixels_7_30, pixels_7_31, pixels_8_0, pixels_8_1, pixels_8_2, pixels_8_3, pixels_8_4, pixels_8_5, pixels_8_6, pixels_8_7, pixels_8_8, pixels_8_9, pixels_8_10, pixels_8_11, pixels_8_12, pixels_8_13, pixels_8_14, pixels_8_15, pixels_8_16, pixels_8_17, pixels_8_18, pixels_8_19, pixels_8_20, pixels_8_21, pixels_8_22, pixels_8_23, pixels_8_24, pixels_8_25, pixels_8_26, pixels_8_27, pixels_8_28, pixels_8_29, pixels_8_30, pixels_8_31, pixels_9_0, pixels_9_1, pixels_9_2, pixels_9_3, pixels_9_4, pixels_9_5, pixels_9_6, pixels_9_7, pixels_9_8, pixels_9_9, pixels_9_10, pixels_9_11, pixels_9_12, pixels_9_13, pixels_9_14, pixels_9_15, pixels_9_16, pixels_9_17, pixels_9_18, pixels_9_19, pixels_9_20, pixels_9_21, pixels_9_22, pixels_9_23, pixels_9_24, pixels_9_25, pixels_9_26, pixels_9_27, pixels_9_28, pixels_9_29, pixels_9_30, pixels_9_31, pixels_10_0, pixels_10_1, pixels_10_2, pixels_10_3, pixels_10_4, pixels_10_5, pixels_10_6, pixels_10_7, pixels_10_8, pixels_10_9, pixels_10_10, pixels_10_11, pixels_10_12, pixels_10_13, pixels_10_14, pixels_10_15, pixels_10_16, pixels_10_17, pixels_10_18, pixels_10_19, pixels_10_20, pixels_10_21, pixels_10_22, pixels_10_23, pixels_10_24, pixels_10_25, pixels_10_26, pixels_10_27, pixels_10_28, pixels_10_29, pixels_10_30, pixels_10_31, pixels_11_0, pixels_11_1, pixels_11_2, pixels_11_3, pixels_11_4, pixels_11_5, pixels_11_6, pixels_11_7, pixels_11_8, pixels_11_9, pixels_11_10, pixels_11_11, pixels_11_12, pixels_11_13, pixels_11_14, pixels_11_15, pixels_11_16, pixels_11_17, pixels_11_18, pixels_11_19, pixels_11_20, pixels_11_21, pixels_11_22, pixels_11_23, pixels_11_24, pixels_11_25, pixels_11_26, pixels_11_27, pixels_11_28, pixels_11_29, pixels_11_30, pixels_11_31, pixels_12_0, pixels_12_1, pixels_12_2, pixels_12_3, pixels_12_4, pixels_12_5, pixels_12_6, pixels_12_7, pixels_12_8, pixels_12_9, pixels_12_10, pixels_12_11, pixels_12_12, pixels_12_13, pixels_12_14, pixels_12_15, pixels_12_16, pixels_12_17, pixels_12_18, pixels_12_19, pixels_12_20, pixels_12_21, pixels_12_22, pixels_12_23, pixels_12_24, pixels_12_25, pixels_12_26, pixels_12_27, pixels_12_28, pixels_12_29, pixels_12_30, pixels_12_31, pixels_13_0, pixels_13_1, pixels_13_2, pixels_13_3, pixels_13_4, pixels_13_5, pixels_13_6, pixels_13_7, pixels_13_8, pixels_13_9, pixels_13_10, pixels_13_11, pixels_13_12, pixels_13_13, pixels_13_14, pixels_13_15, pixels_13_16, pixels_13_17, pixels_13_18, pixels_13_19, pixels_13_20, pixels_13_21, pixels_13_22, pixels_13_23, pixels_13_24, pixels_13_25, pixels_13_26, pixels_13_27, pixels_13_28, pixels_13_29, pixels_13_30, pixels_13_31, pixels_14_0, pixels_14_1, pixels_14_2, pixels_14_3, pixels_14_4, pixels_14_5, pixels_14_6, pixels_14_7, pixels_14_8, pixels_14_9, pixels_14_10, pixels_14_11, pixels_14_12, pixels_14_13, pixels_14_14, pixels_14_15, pixels_14_16, pixels_14_17, pixels_14_18, pixels_14_19, pixels_14_20, pixels_14_21, pixels_14_22, pixels_14_23, pixels_14_24, pixels_14_25, pixels_14_26, pixels_14_27, pixels_14_28, pixels_14_29, pixels_14_30, pixels_14_31, pixels_15_0, pixels_15_1, pixels_15_2, pixels_15_3, pixels_15_4, pixels_15_5, pixels_15_6, pixels_15_7, pixels_15_8, pixels_15_9, pixels_15_10, pixels_15_11, pixels_15_12, pixels_15_13, pixels_15_14, pixels_15_15, pixels_15_16, pixels_15_17, pixels_15_18, pixels_15_19, pixels_15_20, pixels_15_21, pixels_15_22, pixels_15_23, pixels_15_24, pixels_15_25, pixels_15_26, pixels_15_27, pixels_15_28, pixels_15_29, pixels_15_30, pixels_15_31, pixels_16_0, pixels_16_1, pixels_16_2, pixels_16_3, pixels_16_4, pixels_16_5, pixels_16_6, pixels_16_7, pixels_16_8, pixels_16_9, pixels_16_10, pixels_16_11, pixels_16_12, pixels_16_13, pixels_16_14, pixels_16_15, pixels_16_16, pixels_16_17, pixels_16_18, pixels_16_19, pixels_16_20, pixels_16_21, pixels_16_22, pixels_16_23, pixels_16_24, pixels_16_25, pixels_16_26, pixels_16_27, pixels_16_28, pixels_16_29, pixels_16_30, pixels_16_31, pixels_17_0, pixels_17_1, pixels_17_2, pixels_17_3, pixels_17_4, pixels_17_5, pixels_17_6, pixels_17_7, pixels_17_8, pixels_17_9, pixels_17_10, pixels_17_11, pixels_17_12, pixels_17_13, pixels_17_14, pixels_17_15, pixels_17_16, pixels_17_17, pixels_17_18, pixels_17_19, pixels_17_20, pixels_17_21, pixels_17_22, pixels_17_23, pixels_17_24, pixels_17_25, pixels_17_26, pixels_17_27, pixels_17_28, pixels_17_29, pixels_17_30, pixels_17_31, pixels_18_0, pixels_18_1, pixels_18_2, pixels_18_3, pixels_18_4, pixels_18_5, pixels_18_6, pixels_18_7, pixels_18_8, pixels_18_9, pixels_18_10, pixels_18_11, pixels_18_12, pixels_18_13, pixels_18_14, pixels_18_15, pixels_18_16, pixels_18_17, pixels_18_18, pixels_18_19, pixels_18_20, pixels_18_21, pixels_18_22, pixels_18_23, pixels_18_24, pixels_18_25, pixels_18_26, pixels_18_27, pixels_18_28, pixels_18_29, pixels_18_30, pixels_18_31, pixels_19_0, pixels_19_1, pixels_19_2, pixels_19_3, pixels_19_4, pixels_19_5, pixels_19_6, pixels_19_7, pixels_19_8, pixels_19_9, pixels_19_10, pixels_19_11, pixels_19_12, pixels_19_13, pixels_19_14, pixels_19_15, pixels_19_16, pixels_19_17, pixels_19_18, pixels_19_19, pixels_19_20, pixels_19_21, pixels_19_22, pixels_19_23, pixels_19_24, pixels_19_25, pixels_19_26, pixels_19_27, pixels_19_28, pixels_19_29, pixels_19_30, pixels_19_31, pixels_20_0, pixels_20_1, pixels_20_2, pixels_20_3, pixels_20_4, pixels_20_5, pixels_20_6, pixels_20_7, pixels_20_8, pixels_20_9, pixels_20_10, pixels_20_11, pixels_20_12, pixels_20_13, pixels_20_14, pixels_20_15, pixels_20_16, pixels_20_17, pixels_20_18, pixels_20_19, pixels_20_20, pixels_20_21, pixels_20_22, pixels_20_23, pixels_20_24, pixels_20_25, pixels_20_26, pixels_20_27, pixels_20_28, pixels_20_29, pixels_20_30, pixels_20_31, pixels_21_0, pixels_21_1, pixels_21_2, pixels_21_3, pixels_21_4, pixels_21_5, pixels_21_6, pixels_21_7, pixels_21_8, pixels_21_9, pixels_21_10, pixels_21_11, pixels_21_12, pixels_21_13, pixels_21_14, pixels_21_15, pixels_21_16, pixels_21_17, pixels_21_18, pixels_21_19, pixels_21_20, pixels_21_21, pixels_21_22, pixels_21_23, pixels_21_24, pixels_21_25, pixels_21_26, pixels_21_27, pixels_21_28, pixels_21_29, pixels_21_30, pixels_21_31, pixels_22_0, pixels_22_1, pixels_22_2, pixels_22_3, pixels_22_4, pixels_22_5, pixels_22_6, pixels_22_7, pixels_22_8, pixels_22_9, pixels_22_10, pixels_22_11, pixels_22_12, pixels_22_13, pixels_22_14, pixels_22_15, pixels_22_16, pixels_22_17, pixels_22_18, pixels_22_19, pixels_22_20, pixels_22_21, pixels_22_22, pixels_22_23, pixels_22_24, pixels_22_25, pixels_22_26, pixels_22_27, pixels_22_28, pixels_22_29, pixels_22_30, pixels_22_31, 
pixels_23_0, pixels_23_1, pixels_23_2, pixels_23_3, pixels_23_4, pixels_23_5, pixels_23_6, pixels_23_7, pixels_23_8, pixels_23_9, pixels_23_10, pixels_23_11, pixels_23_12, pixels_23_13, pixels_23_14, pixels_23_15, pixels_23_16, pixels_23_17, pixels_23_18, pixels_23_19, pixels_23_20, pixels_23_21, pixels_23_22, pixels_23_23, pixels_23_24, pixels_23_25, pixels_23_26, pixels_23_27, pixels_23_28, pixels_23_29, pixels_23_30, pixels_23_31, pixels_24_0, pixels_24_1, pixels_24_2, pixels_24_3, pixels_24_4, pixels_24_5, pixels_24_6, pixels_24_7, pixels_24_8, pixels_24_9, pixels_24_10, pixels_24_11, pixels_24_12, pixels_24_13, pixels_24_14, pixels_24_15, pixels_24_16, pixels_24_17, pixels_24_18, pixels_24_19, pixels_24_20, pixels_24_21, pixels_24_22, pixels_24_23, pixels_24_24, pixels_24_25, pixels_24_26, pixels_24_27, pixels_24_28, pixels_24_29, pixels_24_30, pixels_24_31, pixels_25_0, pixels_25_1, pixels_25_2, pixels_25_3, pixels_25_4, pixels_25_5, pixels_25_6, pixels_25_7, pixels_25_8, pixels_25_9, pixels_25_10, pixels_25_11, pixels_25_12, pixels_25_13, pixels_25_14, pixels_25_15, pixels_25_16, pixels_25_17, pixels_25_18, pixels_25_19, pixels_25_20, pixels_25_21, pixels_25_22, pixels_25_23, pixels_25_24, pixels_25_25, pixels_25_26, pixels_25_27, pixels_25_28, pixels_25_29, pixels_25_30, pixels_25_31, pixels_26_0, pixels_26_1, pixels_26_2, pixels_26_3, pixels_26_4, pixels_26_5, pixels_26_6, pixels_26_7, pixels_26_8, pixels_26_9, pixels_26_10, pixels_26_11, pixels_26_12, pixels_26_13, pixels_26_14, pixels_26_15, pixels_26_16, pixels_26_17, pixels_26_18, pixels_26_19, pixels_26_20, pixels_26_21, pixels_26_22, pixels_26_23, pixels_26_24, pixels_26_25, pixels_26_26, pixels_26_27, pixels_26_28, pixels_26_29, pixels_26_30, pixels_26_31, pixels_27_0, pixels_27_1, pixels_27_2, pixels_27_3, pixels_27_4, pixels_27_5, pixels_27_6, pixels_27_7, pixels_27_8, pixels_27_9, pixels_27_10, pixels_27_11, pixels_27_12, pixels_27_13, pixels_27_14, pixels_27_15, pixels_27_16, pixels_27_17, pixels_27_18, pixels_27_19, pixels_27_20, pixels_27_21, pixels_27_22, pixels_27_23, pixels_27_24, pixels_27_25, pixels_27_26, pixels_27_27, pixels_27_28, pixels_27_29, pixels_27_30, pixels_27_31, pixels_28_0, pixels_28_1, pixels_28_2, pixels_28_3, pixels_28_4, pixels_28_5, pixels_28_6, pixels_28_7, pixels_28_8, pixels_28_9, pixels_28_10, pixels_28_11, pixels_28_12, pixels_28_13, pixels_28_14, pixels_28_15, pixels_28_16, pixels_28_17, pixels_28_18, pixels_28_19, pixels_28_20, pixels_28_21, pixels_28_22, pixels_28_23, pixels_28_24, pixels_28_25, pixels_28_26, pixels_28_27, pixels_28_28, pixels_28_29, pixels_28_30, pixels_28_31, pixels_29_0, pixels_29_1, pixels_29_2, pixels_29_3, pixels_29_4, pixels_29_5, pixels_29_6, pixels_29_7, pixels_29_8, pixels_29_9, pixels_29_10, pixels_29_11, pixels_29_12, pixels_29_13, pixels_29_14, pixels_29_15, pixels_29_16, pixels_29_17, pixels_29_18, pixels_29_19, pixels_29_20, pixels_29_21, pixels_29_22, pixels_29_23, pixels_29_24, pixels_29_25, pixels_29_26, pixels_29_27, pixels_29_28, pixels_29_29, pixels_29_30, pixels_29_31, pixels_30_0, pixels_30_1, pixels_30_2, pixels_30_3, pixels_30_4, pixels_30_5, pixels_30_6, pixels_30_7, pixels_30_8, pixels_30_9, pixels_30_10, pixels_30_11, pixels_30_12, pixels_30_13, pixels_30_14, pixels_30_15, pixels_30_16, pixels_30_17, pixels_30_18, pixels_30_19, pixels_30_20, pixels_30_21, pixels_30_22, pixels_30_23, pixels_30_24, pixels_30_25, pixels_30_26, pixels_30_27, pixels_30_28, pixels_30_29, pixels_30_30, pixels_30_31, pixels_31_0, pixels_31_1, pixels_31_2, pixels_31_3, pixels_31_4, pixels_31_5, pixels_31_6, pixels_31_7, pixels_31_8, pixels_31_9, pixels_31_10, pixels_31_11, pixels_31_12, pixels_31_13, pixels_31_14, pixels_31_15, pixels_31_16, pixels_31_17, pixels_31_18, pixels_31_19, pixels_31_20, pixels_31_21, pixels_31_22, pixels_31_23, pixels_31_24, pixels_31_25, pixels_31_26, pixels_31_27, pixels_31_28, pixels_31_29, pixels_31_30, pixels_31_31;

wire [(image_size-(kernel_size-kernel_size%2))*(image_size-(kernel_size-kernel_size%2))*word_length*2-1:0] data_out;

assign pixels_0_0 = {data_out[1*word_length*2-1 -: word_length*2]};
assign pixels_1_0 = {data_out[2*word_length*2-1 -: word_length*2]};
assign pixels_2_0 = {data_out[3*word_length*2-1 -: word_length*2]};
assign pixels_3_0 = {data_out[4*word_length*2-1 -: word_length*2]};
assign pixels_4_0 = {data_out[5*word_length*2-1 -: word_length*2]};
assign pixels_5_0 = {data_out[6*word_length*2-1 -: word_length*2]};
assign pixels_6_0 = {data_out[7*word_length*2-1 -: word_length*2]};
assign pixels_7_0 = {data_out[8*word_length*2-1 -: word_length*2]};
assign pixels_8_0 = {data_out[9*word_length*2-1 -: word_length*2]};
assign pixels_9_0 = {data_out[10*word_length*2-1 -: word_length*2]};
assign pixels_10_0 = {data_out[11*word_length*2-1 -: word_length*2]};
assign pixels_11_0 = {data_out[12*word_length*2-1 -: word_length*2]};
assign pixels_12_0 = {data_out[13*word_length*2-1 -: word_length*2]};
assign pixels_13_0 = {data_out[14*word_length*2-1 -: word_length*2]};
assign pixels_14_0 = {data_out[15*word_length*2-1 -: word_length*2]};
assign pixels_15_0 = {data_out[16*word_length*2-1 -: word_length*2]};
assign pixels_16_0 = {data_out[17*word_length*2-1 -: word_length*2]};
assign pixels_17_0 = {data_out[18*word_length*2-1 -: word_length*2]};
assign pixels_18_0 = {data_out[19*word_length*2-1 -: word_length*2]};
assign pixels_19_0 = {data_out[20*word_length*2-1 -: word_length*2]};
assign pixels_20_0 = {data_out[21*word_length*2-1 -: word_length*2]};
assign pixels_21_0 = {data_out[22*word_length*2-1 -: word_length*2]};
assign pixels_22_0 = {data_out[23*word_length*2-1 -: word_length*2]};
assign pixels_23_0 = {data_out[24*word_length*2-1 -: word_length*2]};
assign pixels_24_0 = {data_out[25*word_length*2-1 -: word_length*2]};
assign pixels_25_0 = {data_out[26*word_length*2-1 -: word_length*2]};
assign pixels_26_0 = {data_out[27*word_length*2-1 -: word_length*2]};
assign pixels_27_0 = {data_out[28*word_length*2-1 -: word_length*2]};
assign pixels_28_0 = {data_out[29*word_length*2-1 -: word_length*2]};
assign pixels_29_0 = {data_out[30*word_length*2-1 -: word_length*2]};
assign pixels_30_0 = {data_out[31*word_length*2-1 -: word_length*2]};
assign pixels_31_0 = {data_out[32*word_length*2-1 -: word_length*2]};
assign pixels_0_1 = {data_out[33*word_length*2-1 -: word_length*2]};
assign pixels_1_1 = {data_out[34*word_length*2-1 -: word_length*2]};
assign pixels_2_1 = {data_out[35*word_length*2-1 -: word_length*2]};
assign pixels_3_1 = {data_out[36*word_length*2-1 -: word_length*2]};
assign pixels_4_1 = {data_out[37*word_length*2-1 -: word_length*2]};
assign pixels_5_1 = {data_out[38*word_length*2-1 -: word_length*2]};
assign pixels_6_1 = {data_out[39*word_length*2-1 -: word_length*2]};
assign pixels_7_1 = {data_out[40*word_length*2-1 -: word_length*2]};
assign pixels_8_1 = {data_out[41*word_length*2-1 -: word_length*2]};
assign pixels_9_1 = {data_out[42*word_length*2-1 -: word_length*2]};
assign pixels_10_1 = {data_out[43*word_length*2-1 -: word_length*2]};
assign pixels_11_1 = {data_out[44*word_length*2-1 -: word_length*2]};
assign pixels_12_1 = {data_out[45*word_length*2-1 -: word_length*2]};
assign pixels_13_1 = {data_out[46*word_length*2-1 -: word_length*2]};
assign pixels_14_1 = {data_out[47*word_length*2-1 -: word_length*2]};
assign pixels_15_1 = {data_out[48*word_length*2-1 -: word_length*2]};
assign pixels_16_1 = {data_out[49*word_length*2-1 -: word_length*2]};
assign pixels_17_1 = {data_out[50*word_length*2-1 -: word_length*2]};
assign pixels_18_1 = {data_out[51*word_length*2-1 -: word_length*2]};
assign pixels_19_1 = {data_out[52*word_length*2-1 -: word_length*2]};
assign pixels_20_1 = {data_out[53*word_length*2-1 -: word_length*2]};
assign pixels_21_1 = {data_out[54*word_length*2-1 -: word_length*2]};
assign pixels_22_1 = {data_out[55*word_length*2-1 -: word_length*2]};
assign pixels_23_1 = {data_out[56*word_length*2-1 -: word_length*2]};
assign pixels_24_1 = {data_out[57*word_length*2-1 -: word_length*2]};
assign pixels_25_1 = {data_out[58*word_length*2-1 -: word_length*2]};
assign pixels_26_1 = {data_out[59*word_length*2-1 -: word_length*2]};
assign pixels_27_1 = {data_out[60*word_length*2-1 -: word_length*2]};
assign pixels_28_1 = {data_out[61*word_length*2-1 -: word_length*2]};
assign pixels_29_1 = {data_out[62*word_length*2-1 -: word_length*2]};
assign pixels_30_1 = {data_out[63*word_length*2-1 -: word_length*2]};
assign pixels_31_1 = {data_out[64*word_length*2-1 -: word_length*2]};
assign pixels_0_2 = {data_out[65*word_length*2-1 -: word_length*2]};
assign pixels_1_2 = {data_out[66*word_length*2-1 -: word_length*2]};
assign pixels_2_2 = {data_out[67*word_length*2-1 -: word_length*2]};
assign pixels_3_2 = {data_out[68*word_length*2-1 -: word_length*2]};
assign pixels_4_2 = {data_out[69*word_length*2-1 -: word_length*2]};
assign pixels_5_2 = {data_out[70*word_length*2-1 -: word_length*2]};
assign pixels_6_2 = {data_out[71*word_length*2-1 -: word_length*2]};
assign pixels_7_2 = {data_out[72*word_length*2-1 -: word_length*2]};
assign pixels_8_2 = {data_out[73*word_length*2-1 -: word_length*2]};
assign pixels_9_2 = {data_out[74*word_length*2-1 -: word_length*2]};
assign pixels_10_2 = {data_out[75*word_length*2-1 -: word_length*2]};
assign pixels_11_2 = {data_out[76*word_length*2-1 -: word_length*2]};
assign pixels_12_2 = {data_out[77*word_length*2-1 -: word_length*2]};
assign pixels_13_2 = {data_out[78*word_length*2-1 -: word_length*2]};
assign pixels_14_2 = {data_out[79*word_length*2-1 -: word_length*2]};
assign pixels_15_2 = {data_out[80*word_length*2-1 -: word_length*2]};
assign pixels_16_2 = {data_out[81*word_length*2-1 -: word_length*2]};
assign pixels_17_2 = {data_out[82*word_length*2-1 -: word_length*2]};
assign pixels_18_2 = {data_out[83*word_length*2-1 -: word_length*2]};
assign pixels_19_2 = {data_out[84*word_length*2-1 -: word_length*2]};
assign pixels_20_2 = {data_out[85*word_length*2-1 -: word_length*2]};
assign pixels_21_2 = {data_out[86*word_length*2-1 -: word_length*2]};
assign pixels_22_2 = {data_out[87*word_length*2-1 -: word_length*2]};
assign pixels_23_2 = {data_out[88*word_length*2-1 -: word_length*2]};
assign pixels_24_2 = {data_out[89*word_length*2-1 -: word_length*2]};
assign pixels_25_2 = {data_out[90*word_length*2-1 -: word_length*2]};
assign pixels_26_2 = {data_out[91*word_length*2-1 -: word_length*2]};
assign pixels_27_2 = {data_out[92*word_length*2-1 -: word_length*2]};
assign pixels_28_2 = {data_out[93*word_length*2-1 -: word_length*2]};
assign pixels_29_2 = {data_out[94*word_length*2-1 -: word_length*2]};
assign pixels_30_2 = {data_out[95*word_length*2-1 -: word_length*2]};
assign pixels_31_2 = {data_out[96*word_length*2-1 -: word_length*2]};
assign pixels_0_3 = {data_out[97*word_length*2-1 -: word_length*2]};
assign pixels_1_3 = {data_out[98*word_length*2-1 -: word_length*2]};
assign pixels_2_3 = {data_out[99*word_length*2-1 -: word_length*2]};
assign pixels_3_3 = {data_out[100*word_length*2-1 -: word_length*2]};
assign pixels_4_3 = {data_out[101*word_length*2-1 -: word_length*2]};
assign pixels_5_3 = {data_out[102*word_length*2-1 -: word_length*2]};
assign pixels_6_3 = {data_out[103*word_length*2-1 -: word_length*2]};
assign pixels_7_3 = {data_out[104*word_length*2-1 -: word_length*2]};
assign pixels_8_3 = {data_out[105*word_length*2-1 -: word_length*2]};
assign pixels_9_3 = {data_out[106*word_length*2-1 -: word_length*2]};
assign pixels_10_3 = {data_out[107*word_length*2-1 -: word_length*2]};
assign pixels_11_3 = {data_out[108*word_length*2-1 -: word_length*2]};
assign pixels_12_3 = {data_out[109*word_length*2-1 -: word_length*2]};
assign pixels_13_3 = {data_out[110*word_length*2-1 -: word_length*2]};
assign pixels_14_3 = {data_out[111*word_length*2-1 -: word_length*2]};
assign pixels_15_3 = {data_out[112*word_length*2-1 -: word_length*2]};
assign pixels_16_3 = {data_out[113*word_length*2-1 -: word_length*2]};
assign pixels_17_3 = {data_out[114*word_length*2-1 -: word_length*2]};
assign pixels_18_3 = {data_out[115*word_length*2-1 -: word_length*2]};
assign pixels_19_3 = {data_out[116*word_length*2-1 -: word_length*2]};
assign pixels_20_3 = {data_out[117*word_length*2-1 -: word_length*2]};
assign pixels_21_3 = {data_out[118*word_length*2-1 -: word_length*2]};
assign pixels_22_3 = {data_out[119*word_length*2-1 -: word_length*2]};
assign pixels_23_3 = {data_out[120*word_length*2-1 -: word_length*2]};
assign pixels_24_3 = {data_out[121*word_length*2-1 -: word_length*2]};
assign pixels_25_3 = {data_out[122*word_length*2-1 -: word_length*2]};
assign pixels_26_3 = {data_out[123*word_length*2-1 -: word_length*2]};
assign pixels_27_3 = {data_out[124*word_length*2-1 -: word_length*2]};
assign pixels_28_3 = {data_out[125*word_length*2-1 -: word_length*2]};
assign pixels_29_3 = {data_out[126*word_length*2-1 -: word_length*2]};
assign pixels_30_3 = {data_out[127*word_length*2-1 -: word_length*2]};
assign pixels_31_3 = {data_out[128*word_length*2-1 -: word_length*2]};
assign pixels_0_4 = {data_out[129*word_length*2-1 -: word_length*2]};
assign pixels_1_4 = {data_out[130*word_length*2-1 -: word_length*2]};
assign pixels_2_4 = {data_out[131*word_length*2-1 -: word_length*2]};
assign pixels_3_4 = {data_out[132*word_length*2-1 -: word_length*2]};
assign pixels_4_4 = {data_out[133*word_length*2-1 -: word_length*2]};
assign pixels_5_4 = {data_out[134*word_length*2-1 -: word_length*2]};
assign pixels_6_4 = {data_out[135*word_length*2-1 -: word_length*2]};
assign pixels_7_4 = {data_out[136*word_length*2-1 -: word_length*2]};
assign pixels_8_4 = {data_out[137*word_length*2-1 -: word_length*2]};
assign pixels_9_4 = {data_out[138*word_length*2-1 -: word_length*2]};
assign pixels_10_4 = {data_out[139*word_length*2-1 -: word_length*2]};
assign pixels_11_4 = {data_out[140*word_length*2-1 -: word_length*2]};
assign pixels_12_4 = {data_out[141*word_length*2-1 -: word_length*2]};
assign pixels_13_4 = {data_out[142*word_length*2-1 -: word_length*2]};
assign pixels_14_4 = {data_out[143*word_length*2-1 -: word_length*2]};
assign pixels_15_4 = {data_out[144*word_length*2-1 -: word_length*2]};
assign pixels_16_4 = {data_out[145*word_length*2-1 -: word_length*2]};
assign pixels_17_4 = {data_out[146*word_length*2-1 -: word_length*2]};
assign pixels_18_4 = {data_out[147*word_length*2-1 -: word_length*2]};
assign pixels_19_4 = {data_out[148*word_length*2-1 -: word_length*2]};
assign pixels_20_4 = {data_out[149*word_length*2-1 -: word_length*2]};
assign pixels_21_4 = {data_out[150*word_length*2-1 -: word_length*2]};
assign pixels_22_4 = {data_out[151*word_length*2-1 -: word_length*2]};
assign pixels_23_4 = {data_out[152*word_length*2-1 -: word_length*2]};
assign pixels_24_4 = {data_out[153*word_length*2-1 -: word_length*2]};
assign pixels_25_4 = {data_out[154*word_length*2-1 -: word_length*2]};
assign pixels_26_4 = {data_out[155*word_length*2-1 -: word_length*2]};
assign pixels_27_4 = {data_out[156*word_length*2-1 -: word_length*2]};
assign pixels_28_4 = {data_out[157*word_length*2-1 -: word_length*2]};
assign pixels_29_4 = {data_out[158*word_length*2-1 -: word_length*2]};
assign pixels_30_4 = {data_out[159*word_length*2-1 -: word_length*2]};
assign pixels_31_4 = {data_out[160*word_length*2-1 -: word_length*2]};
assign pixels_0_5 = {data_out[161*word_length*2-1 -: word_length*2]};
assign pixels_1_5 = {data_out[162*word_length*2-1 -: word_length*2]};
assign pixels_2_5 = {data_out[163*word_length*2-1 -: word_length*2]};
assign pixels_3_5 = {data_out[164*word_length*2-1 -: word_length*2]};
assign pixels_4_5 = {data_out[165*word_length*2-1 -: word_length*2]};
assign pixels_5_5 = {data_out[166*word_length*2-1 -: word_length*2]};
assign pixels_6_5 = {data_out[167*word_length*2-1 -: word_length*2]};
assign pixels_7_5 = {data_out[168*word_length*2-1 -: word_length*2]};
assign pixels_8_5 = {data_out[169*word_length*2-1 -: word_length*2]};
assign pixels_9_5 = {data_out[170*word_length*2-1 -: word_length*2]};
assign pixels_10_5 = {data_out[171*word_length*2-1 -: word_length*2]};
assign pixels_11_5 = {data_out[172*word_length*2-1 -: word_length*2]};
assign pixels_12_5 = {data_out[173*word_length*2-1 -: word_length*2]};
assign pixels_13_5 = {data_out[174*word_length*2-1 -: word_length*2]};
assign pixels_14_5 = {data_out[175*word_length*2-1 -: word_length*2]};
assign pixels_15_5 = {data_out[176*word_length*2-1 -: word_length*2]};
assign pixels_16_5 = {data_out[177*word_length*2-1 -: word_length*2]};
assign pixels_17_5 = {data_out[178*word_length*2-1 -: word_length*2]};
assign pixels_18_5 = {data_out[179*word_length*2-1 -: word_length*2]};
assign pixels_19_5 = {data_out[180*word_length*2-1 -: word_length*2]};
assign pixels_20_5 = {data_out[181*word_length*2-1 -: word_length*2]};
assign pixels_21_5 = {data_out[182*word_length*2-1 -: word_length*2]};
assign pixels_22_5 = {data_out[183*word_length*2-1 -: word_length*2]};
assign pixels_23_5 = {data_out[184*word_length*2-1 -: word_length*2]};
assign pixels_24_5 = {data_out[185*word_length*2-1 -: word_length*2]};
assign pixels_25_5 = {data_out[186*word_length*2-1 -: word_length*2]};
assign pixels_26_5 = {data_out[187*word_length*2-1 -: word_length*2]};
assign pixels_27_5 = {data_out[188*word_length*2-1 -: word_length*2]};
assign pixels_28_5 = {data_out[189*word_length*2-1 -: word_length*2]};
assign pixels_29_5 = {data_out[190*word_length*2-1 -: word_length*2]};
assign pixels_30_5 = {data_out[191*word_length*2-1 -: word_length*2]};
assign pixels_31_5 = {data_out[192*word_length*2-1 -: word_length*2]};
assign pixels_0_6 = {data_out[193*word_length*2-1 -: word_length*2]};
assign pixels_1_6 = {data_out[194*word_length*2-1 -: word_length*2]};
assign pixels_2_6 = {data_out[195*word_length*2-1 -: word_length*2]};
assign pixels_3_6 = {data_out[196*word_length*2-1 -: word_length*2]};
assign pixels_4_6 = {data_out[197*word_length*2-1 -: word_length*2]};
assign pixels_5_6 = {data_out[198*word_length*2-1 -: word_length*2]};
assign pixels_6_6 = {data_out[199*word_length*2-1 -: word_length*2]};
assign pixels_7_6 = {data_out[200*word_length*2-1 -: word_length*2]};
assign pixels_8_6 = {data_out[201*word_length*2-1 -: word_length*2]};
assign pixels_9_6 = {data_out[202*word_length*2-1 -: word_length*2]};
assign pixels_10_6 = {data_out[203*word_length*2-1 -: word_length*2]};
assign pixels_11_6 = {data_out[204*word_length*2-1 -: word_length*2]};
assign pixels_12_6 = {data_out[205*word_length*2-1 -: word_length*2]};
assign pixels_13_6 = {data_out[206*word_length*2-1 -: word_length*2]};
assign pixels_14_6 = {data_out[207*word_length*2-1 -: word_length*2]};
assign pixels_15_6 = {data_out[208*word_length*2-1 -: word_length*2]};
assign pixels_16_6 = {data_out[209*word_length*2-1 -: word_length*2]};
assign pixels_17_6 = {data_out[210*word_length*2-1 -: word_length*2]};
assign pixels_18_6 = {data_out[211*word_length*2-1 -: word_length*2]};
assign pixels_19_6 = {data_out[212*word_length*2-1 -: word_length*2]};
assign pixels_20_6 = {data_out[213*word_length*2-1 -: word_length*2]};
assign pixels_21_6 = {data_out[214*word_length*2-1 -: word_length*2]};
assign pixels_22_6 = {data_out[215*word_length*2-1 -: word_length*2]};
assign pixels_23_6 = {data_out[216*word_length*2-1 -: word_length*2]};
assign pixels_24_6 = {data_out[217*word_length*2-1 -: word_length*2]};
assign pixels_25_6 = {data_out[218*word_length*2-1 -: word_length*2]};
assign pixels_26_6 = {data_out[219*word_length*2-1 -: word_length*2]};
assign pixels_27_6 = {data_out[220*word_length*2-1 -: word_length*2]};
assign pixels_28_6 = {data_out[221*word_length*2-1 -: word_length*2]};
assign pixels_29_6 = {data_out[222*word_length*2-1 -: word_length*2]};
assign pixels_30_6 = {data_out[223*word_length*2-1 -: word_length*2]};
assign pixels_31_6 = {data_out[224*word_length*2-1 -: word_length*2]};
assign pixels_0_7 = {data_out[225*word_length*2-1 -: word_length*2]};
assign pixels_1_7 = {data_out[226*word_length*2-1 -: word_length*2]};
assign pixels_2_7 = {data_out[227*word_length*2-1 -: word_length*2]};
assign pixels_3_7 = {data_out[228*word_length*2-1 -: word_length*2]};
assign pixels_4_7 = {data_out[229*word_length*2-1 -: word_length*2]};
assign pixels_5_7 = {data_out[230*word_length*2-1 -: word_length*2]};
assign pixels_6_7 = {data_out[231*word_length*2-1 -: word_length*2]};
assign pixels_7_7 = {data_out[232*word_length*2-1 -: word_length*2]};
assign pixels_8_7 = {data_out[233*word_length*2-1 -: word_length*2]};
assign pixels_9_7 = {data_out[234*word_length*2-1 -: word_length*2]};
assign pixels_10_7 = {data_out[235*word_length*2-1 -: word_length*2]};
assign pixels_11_7 = {data_out[236*word_length*2-1 -: word_length*2]};
assign pixels_12_7 = {data_out[237*word_length*2-1 -: word_length*2]};
assign pixels_13_7 = {data_out[238*word_length*2-1 -: word_length*2]};
assign pixels_14_7 = {data_out[239*word_length*2-1 -: word_length*2]};
assign pixels_15_7 = {data_out[240*word_length*2-1 -: word_length*2]};
assign pixels_16_7 = {data_out[241*word_length*2-1 -: word_length*2]};
assign pixels_17_7 = {data_out[242*word_length*2-1 -: word_length*2]};
assign pixels_18_7 = {data_out[243*word_length*2-1 -: word_length*2]};
assign pixels_19_7 = {data_out[244*word_length*2-1 -: word_length*2]};
assign pixels_20_7 = {data_out[245*word_length*2-1 -: word_length*2]};
assign pixels_21_7 = {data_out[246*word_length*2-1 -: word_length*2]};
assign pixels_22_7 = {data_out[247*word_length*2-1 -: word_length*2]};
assign pixels_23_7 = {data_out[248*word_length*2-1 -: word_length*2]};
assign pixels_24_7 = {data_out[249*word_length*2-1 -: word_length*2]};
assign pixels_25_7 = {data_out[250*word_length*2-1 -: word_length*2]};
assign pixels_26_7 = {data_out[251*word_length*2-1 -: word_length*2]};
assign pixels_27_7 = {data_out[252*word_length*2-1 -: word_length*2]};
assign pixels_28_7 = {data_out[253*word_length*2-1 -: word_length*2]};
assign pixels_29_7 = {data_out[254*word_length*2-1 -: word_length*2]};
assign pixels_30_7 = {data_out[255*word_length*2-1 -: word_length*2]};
assign pixels_31_7 = {data_out[256*word_length*2-1 -: word_length*2]};
assign pixels_0_8 = {data_out[257*word_length*2-1 -: word_length*2]};
assign pixels_1_8 = {data_out[258*word_length*2-1 -: word_length*2]};
assign pixels_2_8 = {data_out[259*word_length*2-1 -: word_length*2]};
assign pixels_3_8 = {data_out[260*word_length*2-1 -: word_length*2]};
assign pixels_4_8 = {data_out[261*word_length*2-1 -: word_length*2]};
assign pixels_5_8 = {data_out[262*word_length*2-1 -: word_length*2]};
assign pixels_6_8 = {data_out[263*word_length*2-1 -: word_length*2]};
assign pixels_7_8 = {data_out[264*word_length*2-1 -: word_length*2]};
assign pixels_8_8 = {data_out[265*word_length*2-1 -: word_length*2]};
assign pixels_9_8 = {data_out[266*word_length*2-1 -: word_length*2]};
assign pixels_10_8 = {data_out[267*word_length*2-1 -: word_length*2]};
assign pixels_11_8 = {data_out[268*word_length*2-1 -: word_length*2]};
assign pixels_12_8 = {data_out[269*word_length*2-1 -: word_length*2]};
assign pixels_13_8 = {data_out[270*word_length*2-1 -: word_length*2]};
assign pixels_14_8 = {data_out[271*word_length*2-1 -: word_length*2]};
assign pixels_15_8 = {data_out[272*word_length*2-1 -: word_length*2]};
assign pixels_16_8 = {data_out[273*word_length*2-1 -: word_length*2]};
assign pixels_17_8 = {data_out[274*word_length*2-1 -: word_length*2]};
assign pixels_18_8 = {data_out[275*word_length*2-1 -: word_length*2]};
assign pixels_19_8 = {data_out[276*word_length*2-1 -: word_length*2]};
assign pixels_20_8 = {data_out[277*word_length*2-1 -: word_length*2]};
assign pixels_21_8 = {data_out[278*word_length*2-1 -: word_length*2]};
assign pixels_22_8 = {data_out[279*word_length*2-1 -: word_length*2]};
assign pixels_23_8 = {data_out[280*word_length*2-1 -: word_length*2]};
assign pixels_24_8 = {data_out[281*word_length*2-1 -: word_length*2]};
assign pixels_25_8 = {data_out[282*word_length*2-1 -: word_length*2]};
assign pixels_26_8 = {data_out[283*word_length*2-1 -: word_length*2]};
assign pixels_27_8 = {data_out[284*word_length*2-1 -: word_length*2]};
assign pixels_28_8 = {data_out[285*word_length*2-1 -: word_length*2]};
assign pixels_29_8 = {data_out[286*word_length*2-1 -: word_length*2]};
assign pixels_30_8 = {data_out[287*word_length*2-1 -: word_length*2]};
assign pixels_31_8 = {data_out[288*word_length*2-1 -: word_length*2]};
assign pixels_0_9 = {data_out[289*word_length*2-1 -: word_length*2]};
assign pixels_1_9 = {data_out[290*word_length*2-1 -: word_length*2]};
assign pixels_2_9 = {data_out[291*word_length*2-1 -: word_length*2]};
assign pixels_3_9 = {data_out[292*word_length*2-1 -: word_length*2]};
assign pixels_4_9 = {data_out[293*word_length*2-1 -: word_length*2]};
assign pixels_5_9 = {data_out[294*word_length*2-1 -: word_length*2]};
assign pixels_6_9 = {data_out[295*word_length*2-1 -: word_length*2]};
assign pixels_7_9 = {data_out[296*word_length*2-1 -: word_length*2]};
assign pixels_8_9 = {data_out[297*word_length*2-1 -: word_length*2]};
assign pixels_9_9 = {data_out[298*word_length*2-1 -: word_length*2]};
assign pixels_10_9 = {data_out[299*word_length*2-1 -: word_length*2]};
assign pixels_11_9 = {data_out[300*word_length*2-1 -: word_length*2]};
assign pixels_12_9 = {data_out[301*word_length*2-1 -: word_length*2]};
assign pixels_13_9 = {data_out[302*word_length*2-1 -: word_length*2]};
assign pixels_14_9 = {data_out[303*word_length*2-1 -: word_length*2]};
assign pixels_15_9 = {data_out[304*word_length*2-1 -: word_length*2]};
assign pixels_16_9 = {data_out[305*word_length*2-1 -: word_length*2]};
assign pixels_17_9 = {data_out[306*word_length*2-1 -: word_length*2]};
assign pixels_18_9 = {data_out[307*word_length*2-1 -: word_length*2]};
assign pixels_19_9 = {data_out[308*word_length*2-1 -: word_length*2]};
assign pixels_20_9 = {data_out[309*word_length*2-1 -: word_length*2]};
assign pixels_21_9 = {data_out[310*word_length*2-1 -: word_length*2]};
assign pixels_22_9 = {data_out[311*word_length*2-1 -: word_length*2]};
assign pixels_23_9 = {data_out[312*word_length*2-1 -: word_length*2]};
assign pixels_24_9 = {data_out[313*word_length*2-1 -: word_length*2]};
assign pixels_25_9 = {data_out[314*word_length*2-1 -: word_length*2]};
assign pixels_26_9 = {data_out[315*word_length*2-1 -: word_length*2]};
assign pixels_27_9 = {data_out[316*word_length*2-1 -: word_length*2]};
assign pixels_28_9 = {data_out[317*word_length*2-1 -: word_length*2]};
assign pixels_29_9 = {data_out[318*word_length*2-1 -: word_length*2]};
assign pixels_30_9 = {data_out[319*word_length*2-1 -: word_length*2]};
assign pixels_31_9 = {data_out[320*word_length*2-1 -: word_length*2]};
assign pixels_0_10 = {data_out[321*word_length*2-1 -: word_length*2]};
assign pixels_1_10 = {data_out[322*word_length*2-1 -: word_length*2]};
assign pixels_2_10 = {data_out[323*word_length*2-1 -: word_length*2]};
assign pixels_3_10 = {data_out[324*word_length*2-1 -: word_length*2]};
assign pixels_4_10 = {data_out[325*word_length*2-1 -: word_length*2]};
assign pixels_5_10 = {data_out[326*word_length*2-1 -: word_length*2]};
assign pixels_6_10 = {data_out[327*word_length*2-1 -: word_length*2]};
assign pixels_7_10 = {data_out[328*word_length*2-1 -: word_length*2]};
assign pixels_8_10 = {data_out[329*word_length*2-1 -: word_length*2]};
assign pixels_9_10 = {data_out[330*word_length*2-1 -: word_length*2]};
assign pixels_10_10 = {data_out[331*word_length*2-1 -: word_length*2]};
assign pixels_11_10 = {data_out[332*word_length*2-1 -: word_length*2]};
assign pixels_12_10 = {data_out[333*word_length*2-1 -: word_length*2]};
assign pixels_13_10 = {data_out[334*word_length*2-1 -: word_length*2]};
assign pixels_14_10 = {data_out[335*word_length*2-1 -: word_length*2]};
assign pixels_15_10 = {data_out[336*word_length*2-1 -: word_length*2]};
assign pixels_16_10 = {data_out[337*word_length*2-1 -: word_length*2]};
assign pixels_17_10 = {data_out[338*word_length*2-1 -: word_length*2]};
assign pixels_18_10 = {data_out[339*word_length*2-1 -: word_length*2]};
assign pixels_19_10 = {data_out[340*word_length*2-1 -: word_length*2]};
assign pixels_20_10 = {data_out[341*word_length*2-1 -: word_length*2]};
assign pixels_21_10 = {data_out[342*word_length*2-1 -: word_length*2]};
assign pixels_22_10 = {data_out[343*word_length*2-1 -: word_length*2]};
assign pixels_23_10 = {data_out[344*word_length*2-1 -: word_length*2]};
assign pixels_24_10 = {data_out[345*word_length*2-1 -: word_length*2]};
assign pixels_25_10 = {data_out[346*word_length*2-1 -: word_length*2]};
assign pixels_26_10 = {data_out[347*word_length*2-1 -: word_length*2]};
assign pixels_27_10 = {data_out[348*word_length*2-1 -: word_length*2]};
assign pixels_28_10 = {data_out[349*word_length*2-1 -: word_length*2]};
assign pixels_29_10 = {data_out[350*word_length*2-1 -: word_length*2]};
assign pixels_30_10 = {data_out[351*word_length*2-1 -: word_length*2]};
assign pixels_31_10 = {data_out[352*word_length*2-1 -: word_length*2]};
assign pixels_0_11 = {data_out[353*word_length*2-1 -: word_length*2]};
assign pixels_1_11 = {data_out[354*word_length*2-1 -: word_length*2]};
assign pixels_2_11 = {data_out[355*word_length*2-1 -: word_length*2]};
assign pixels_3_11 = {data_out[356*word_length*2-1 -: word_length*2]};
assign pixels_4_11 = {data_out[357*word_length*2-1 -: word_length*2]};
assign pixels_5_11 = {data_out[358*word_length*2-1 -: word_length*2]};
assign pixels_6_11 = {data_out[359*word_length*2-1 -: word_length*2]};
assign pixels_7_11 = {data_out[360*word_length*2-1 -: word_length*2]};
assign pixels_8_11 = {data_out[361*word_length*2-1 -: word_length*2]};
assign pixels_9_11 = {data_out[362*word_length*2-1 -: word_length*2]};
assign pixels_10_11 = {data_out[363*word_length*2-1 -: word_length*2]};
assign pixels_11_11 = {data_out[364*word_length*2-1 -: word_length*2]};
assign pixels_12_11 = {data_out[365*word_length*2-1 -: word_length*2]};
assign pixels_13_11 = {data_out[366*word_length*2-1 -: word_length*2]};
assign pixels_14_11 = {data_out[367*word_length*2-1 -: word_length*2]};
assign pixels_15_11 = {data_out[368*word_length*2-1 -: word_length*2]};
assign pixels_16_11 = {data_out[369*word_length*2-1 -: word_length*2]};
assign pixels_17_11 = {data_out[370*word_length*2-1 -: word_length*2]};
assign pixels_18_11 = {data_out[371*word_length*2-1 -: word_length*2]};
assign pixels_19_11 = {data_out[372*word_length*2-1 -: word_length*2]};
assign pixels_20_11 = {data_out[373*word_length*2-1 -: word_length*2]};
assign pixels_21_11 = {data_out[374*word_length*2-1 -: word_length*2]};
assign pixels_22_11 = {data_out[375*word_length*2-1 -: word_length*2]};
assign pixels_23_11 = {data_out[376*word_length*2-1 -: word_length*2]};
assign pixels_24_11 = {data_out[377*word_length*2-1 -: word_length*2]};
assign pixels_25_11 = {data_out[378*word_length*2-1 -: word_length*2]};
assign pixels_26_11 = {data_out[379*word_length*2-1 -: word_length*2]};
assign pixels_27_11 = {data_out[380*word_length*2-1 -: word_length*2]};
assign pixels_28_11 = {data_out[381*word_length*2-1 -: word_length*2]};
assign pixels_29_11 = {data_out[382*word_length*2-1 -: word_length*2]};
assign pixels_30_11 = {data_out[383*word_length*2-1 -: word_length*2]};
assign pixels_31_11 = {data_out[384*word_length*2-1 -: word_length*2]};
assign pixels_0_12 = {data_out[385*word_length*2-1 -: word_length*2]};
assign pixels_1_12 = {data_out[386*word_length*2-1 -: word_length*2]};
assign pixels_2_12 = {data_out[387*word_length*2-1 -: word_length*2]};
assign pixels_3_12 = {data_out[388*word_length*2-1 -: word_length*2]};
assign pixels_4_12 = {data_out[389*word_length*2-1 -: word_length*2]};
assign pixels_5_12 = {data_out[390*word_length*2-1 -: word_length*2]};
assign pixels_6_12 = {data_out[391*word_length*2-1 -: word_length*2]};
assign pixels_7_12 = {data_out[392*word_length*2-1 -: word_length*2]};
assign pixels_8_12 = {data_out[393*word_length*2-1 -: word_length*2]};
assign pixels_9_12 = {data_out[394*word_length*2-1 -: word_length*2]};
assign pixels_10_12 = {data_out[395*word_length*2-1 -: word_length*2]};
assign pixels_11_12 = {data_out[396*word_length*2-1 -: word_length*2]};
assign pixels_12_12 = {data_out[397*word_length*2-1 -: word_length*2]};
assign pixels_13_12 = {data_out[398*word_length*2-1 -: word_length*2]};
assign pixels_14_12 = {data_out[399*word_length*2-1 -: word_length*2]};
assign pixels_15_12 = {data_out[400*word_length*2-1 -: word_length*2]};
assign pixels_16_12 = {data_out[401*word_length*2-1 -: word_length*2]};
assign pixels_17_12 = {data_out[402*word_length*2-1 -: word_length*2]};
assign pixels_18_12 = {data_out[403*word_length*2-1 -: word_length*2]};
assign pixels_19_12 = {data_out[404*word_length*2-1 -: word_length*2]};
assign pixels_20_12 = {data_out[405*word_length*2-1 -: word_length*2]};
assign pixels_21_12 = {data_out[406*word_length*2-1 -: word_length*2]};
assign pixels_22_12 = {data_out[407*word_length*2-1 -: word_length*2]};
assign pixels_23_12 = {data_out[408*word_length*2-1 -: word_length*2]};
assign pixels_24_12 = {data_out[409*word_length*2-1 -: word_length*2]};
assign pixels_25_12 = {data_out[410*word_length*2-1 -: word_length*2]};
assign pixels_26_12 = {data_out[411*word_length*2-1 -: word_length*2]};
assign pixels_27_12 = {data_out[412*word_length*2-1 -: word_length*2]};
assign pixels_28_12 = {data_out[413*word_length*2-1 -: word_length*2]};
assign pixels_29_12 = {data_out[414*word_length*2-1 -: word_length*2]};
assign pixels_30_12 = {data_out[415*word_length*2-1 -: word_length*2]};
assign pixels_31_12 = {data_out[416*word_length*2-1 -: word_length*2]};
assign pixels_0_13 = {data_out[417*word_length*2-1 -: word_length*2]};
assign pixels_1_13 = {data_out[418*word_length*2-1 -: word_length*2]};
assign pixels_2_13 = {data_out[419*word_length*2-1 -: word_length*2]};
assign pixels_3_13 = {data_out[420*word_length*2-1 -: word_length*2]};
assign pixels_4_13 = {data_out[421*word_length*2-1 -: word_length*2]};
assign pixels_5_13 = {data_out[422*word_length*2-1 -: word_length*2]};
assign pixels_6_13 = {data_out[423*word_length*2-1 -: word_length*2]};
assign pixels_7_13 = {data_out[424*word_length*2-1 -: word_length*2]};
assign pixels_8_13 = {data_out[425*word_length*2-1 -: word_length*2]};
assign pixels_9_13 = {data_out[426*word_length*2-1 -: word_length*2]};
assign pixels_10_13 = {data_out[427*word_length*2-1 -: word_length*2]};
assign pixels_11_13 = {data_out[428*word_length*2-1 -: word_length*2]};
assign pixels_12_13 = {data_out[429*word_length*2-1 -: word_length*2]};
assign pixels_13_13 = {data_out[430*word_length*2-1 -: word_length*2]};
assign pixels_14_13 = {data_out[431*word_length*2-1 -: word_length*2]};
assign pixels_15_13 = {data_out[432*word_length*2-1 -: word_length*2]};
assign pixels_16_13 = {data_out[433*word_length*2-1 -: word_length*2]};
assign pixels_17_13 = {data_out[434*word_length*2-1 -: word_length*2]};
assign pixels_18_13 = {data_out[435*word_length*2-1 -: word_length*2]};
assign pixels_19_13 = {data_out[436*word_length*2-1 -: word_length*2]};
assign pixels_20_13 = {data_out[437*word_length*2-1 -: word_length*2]};
assign pixels_21_13 = {data_out[438*word_length*2-1 -: word_length*2]};
assign pixels_22_13 = {data_out[439*word_length*2-1 -: word_length*2]};
assign pixels_23_13 = {data_out[440*word_length*2-1 -: word_length*2]};
assign pixels_24_13 = {data_out[441*word_length*2-1 -: word_length*2]};
assign pixels_25_13 = {data_out[442*word_length*2-1 -: word_length*2]};
assign pixels_26_13 = {data_out[443*word_length*2-1 -: word_length*2]};
assign pixels_27_13 = {data_out[444*word_length*2-1 -: word_length*2]};
assign pixels_28_13 = {data_out[445*word_length*2-1 -: word_length*2]};
assign pixels_29_13 = {data_out[446*word_length*2-1 -: word_length*2]};
assign pixels_30_13 = {data_out[447*word_length*2-1 -: word_length*2]};
assign pixels_31_13 = {data_out[448*word_length*2-1 -: word_length*2]};
assign pixels_0_14 = {data_out[449*word_length*2-1 -: word_length*2]};
assign pixels_1_14 = {data_out[450*word_length*2-1 -: word_length*2]};
assign pixels_2_14 = {data_out[451*word_length*2-1 -: word_length*2]};
assign pixels_3_14 = {data_out[452*word_length*2-1 -: word_length*2]};
assign pixels_4_14 = {data_out[453*word_length*2-1 -: word_length*2]};
assign pixels_5_14 = {data_out[454*word_length*2-1 -: word_length*2]};
assign pixels_6_14 = {data_out[455*word_length*2-1 -: word_length*2]};
assign pixels_7_14 = {data_out[456*word_length*2-1 -: word_length*2]};
assign pixels_8_14 = {data_out[457*word_length*2-1 -: word_length*2]};
assign pixels_9_14 = {data_out[458*word_length*2-1 -: word_length*2]};
assign pixels_10_14 = {data_out[459*word_length*2-1 -: word_length*2]};
assign pixels_11_14 = {data_out[460*word_length*2-1 -: word_length*2]};
assign pixels_12_14 = {data_out[461*word_length*2-1 -: word_length*2]};
assign pixels_13_14 = {data_out[462*word_length*2-1 -: word_length*2]};
assign pixels_14_14 = {data_out[463*word_length*2-1 -: word_length*2]};
assign pixels_15_14 = {data_out[464*word_length*2-1 -: word_length*2]};
assign pixels_16_14 = {data_out[465*word_length*2-1 -: word_length*2]};
assign pixels_17_14 = {data_out[466*word_length*2-1 -: word_length*2]};
assign pixels_18_14 = {data_out[467*word_length*2-1 -: word_length*2]};
assign pixels_19_14 = {data_out[468*word_length*2-1 -: word_length*2]};
assign pixels_20_14 = {data_out[469*word_length*2-1 -: word_length*2]};
assign pixels_21_14 = {data_out[470*word_length*2-1 -: word_length*2]};
assign pixels_22_14 = {data_out[471*word_length*2-1 -: word_length*2]};
assign pixels_23_14 = {data_out[472*word_length*2-1 -: word_length*2]};
assign pixels_24_14 = {data_out[473*word_length*2-1 -: word_length*2]};
assign pixels_25_14 = {data_out[474*word_length*2-1 -: word_length*2]};
assign pixels_26_14 = {data_out[475*word_length*2-1 -: word_length*2]};
assign pixels_27_14 = {data_out[476*word_length*2-1 -: word_length*2]};
assign pixels_28_14 = {data_out[477*word_length*2-1 -: word_length*2]};
assign pixels_29_14 = {data_out[478*word_length*2-1 -: word_length*2]};
assign pixels_30_14 = {data_out[479*word_length*2-1 -: word_length*2]};
assign pixels_31_14 = {data_out[480*word_length*2-1 -: word_length*2]};
assign pixels_0_15 = {data_out[481*word_length*2-1 -: word_length*2]};
assign pixels_1_15 = {data_out[482*word_length*2-1 -: word_length*2]};
assign pixels_2_15 = {data_out[483*word_length*2-1 -: word_length*2]};
assign pixels_3_15 = {data_out[484*word_length*2-1 -: word_length*2]};
assign pixels_4_15 = {data_out[485*word_length*2-1 -: word_length*2]};
assign pixels_5_15 = {data_out[486*word_length*2-1 -: word_length*2]};
assign pixels_6_15 = {data_out[487*word_length*2-1 -: word_length*2]};
assign pixels_7_15 = {data_out[488*word_length*2-1 -: word_length*2]};
assign pixels_8_15 = {data_out[489*word_length*2-1 -: word_length*2]};
assign pixels_9_15 = {data_out[490*word_length*2-1 -: word_length*2]};
assign pixels_10_15 = {data_out[491*word_length*2-1 -: word_length*2]};
assign pixels_11_15 = {data_out[492*word_length*2-1 -: word_length*2]};
assign pixels_12_15 = {data_out[493*word_length*2-1 -: word_length*2]};
assign pixels_13_15 = {data_out[494*word_length*2-1 -: word_length*2]};
assign pixels_14_15 = {data_out[495*word_length*2-1 -: word_length*2]};
assign pixels_15_15 = {data_out[496*word_length*2-1 -: word_length*2]};
assign pixels_16_15 = {data_out[497*word_length*2-1 -: word_length*2]};
assign pixels_17_15 = {data_out[498*word_length*2-1 -: word_length*2]};
assign pixels_18_15 = {data_out[499*word_length*2-1 -: word_length*2]};
assign pixels_19_15 = {data_out[500*word_length*2-1 -: word_length*2]};
assign pixels_20_15 = {data_out[501*word_length*2-1 -: word_length*2]};
assign pixels_21_15 = {data_out[502*word_length*2-1 -: word_length*2]};
assign pixels_22_15 = {data_out[503*word_length*2-1 -: word_length*2]};
assign pixels_23_15 = {data_out[504*word_length*2-1 -: word_length*2]};
assign pixels_24_15 = {data_out[505*word_length*2-1 -: word_length*2]};
assign pixels_25_15 = {data_out[506*word_length*2-1 -: word_length*2]};
assign pixels_26_15 = {data_out[507*word_length*2-1 -: word_length*2]};
assign pixels_27_15 = {data_out[508*word_length*2-1 -: word_length*2]};
assign pixels_28_15 = {data_out[509*word_length*2-1 -: word_length*2]};
assign pixels_29_15 = {data_out[510*word_length*2-1 -: word_length*2]};
assign pixels_30_15 = {data_out[511*word_length*2-1 -: word_length*2]};
assign pixels_31_15 = {data_out[512*word_length*2-1 -: word_length*2]};
assign pixels_0_16 = {data_out[513*word_length*2-1 -: word_length*2]};
assign pixels_1_16 = {data_out[514*word_length*2-1 -: word_length*2]};
assign pixels_2_16 = {data_out[515*word_length*2-1 -: word_length*2]};
assign pixels_3_16 = {data_out[516*word_length*2-1 -: word_length*2]};
assign pixels_4_16 = {data_out[517*word_length*2-1 -: word_length*2]};
assign pixels_5_16 = {data_out[518*word_length*2-1 -: word_length*2]};
assign pixels_6_16 = {data_out[519*word_length*2-1 -: word_length*2]};
assign pixels_7_16 = {data_out[520*word_length*2-1 -: word_length*2]};
assign pixels_8_16 = {data_out[521*word_length*2-1 -: word_length*2]};
assign pixels_9_16 = {data_out[522*word_length*2-1 -: word_length*2]};
assign pixels_10_16 = {data_out[523*word_length*2-1 -: word_length*2]};
assign pixels_11_16 = {data_out[524*word_length*2-1 -: word_length*2]};
assign pixels_12_16 = {data_out[525*word_length*2-1 -: word_length*2]};
assign pixels_13_16 = {data_out[526*word_length*2-1 -: word_length*2]};
assign pixels_14_16 = {data_out[527*word_length*2-1 -: word_length*2]};
assign pixels_15_16 = {data_out[528*word_length*2-1 -: word_length*2]};
assign pixels_16_16 = {data_out[529*word_length*2-1 -: word_length*2]};
assign pixels_17_16 = {data_out[530*word_length*2-1 -: word_length*2]};
assign pixels_18_16 = {data_out[531*word_length*2-1 -: word_length*2]};
assign pixels_19_16 = {data_out[532*word_length*2-1 -: word_length*2]};
assign pixels_20_16 = {data_out[533*word_length*2-1 -: word_length*2]};
assign pixels_21_16 = {data_out[534*word_length*2-1 -: word_length*2]};
assign pixels_22_16 = {data_out[535*word_length*2-1 -: word_length*2]};
assign pixels_23_16 = {data_out[536*word_length*2-1 -: word_length*2]};
assign pixels_24_16 = {data_out[537*word_length*2-1 -: word_length*2]};
assign pixels_25_16 = {data_out[538*word_length*2-1 -: word_length*2]};
assign pixels_26_16 = {data_out[539*word_length*2-1 -: word_length*2]};
assign pixels_27_16 = {data_out[540*word_length*2-1 -: word_length*2]};
assign pixels_28_16 = {data_out[541*word_length*2-1 -: word_length*2]};
assign pixels_29_16 = {data_out[542*word_length*2-1 -: word_length*2]};
assign pixels_30_16 = {data_out[543*word_length*2-1 -: word_length*2]};
assign pixels_31_16 = {data_out[544*word_length*2-1 -: word_length*2]};
assign pixels_0_17 = {data_out[545*word_length*2-1 -: word_length*2]};
assign pixels_1_17 = {data_out[546*word_length*2-1 -: word_length*2]};
assign pixels_2_17 = {data_out[547*word_length*2-1 -: word_length*2]};
assign pixels_3_17 = {data_out[548*word_length*2-1 -: word_length*2]};
assign pixels_4_17 = {data_out[549*word_length*2-1 -: word_length*2]};
assign pixels_5_17 = {data_out[550*word_length*2-1 -: word_length*2]};
assign pixels_6_17 = {data_out[551*word_length*2-1 -: word_length*2]};
assign pixels_7_17 = {data_out[552*word_length*2-1 -: word_length*2]};
assign pixels_8_17 = {data_out[553*word_length*2-1 -: word_length*2]};
assign pixels_9_17 = {data_out[554*word_length*2-1 -: word_length*2]};
assign pixels_10_17 = {data_out[555*word_length*2-1 -: word_length*2]};
assign pixels_11_17 = {data_out[556*word_length*2-1 -: word_length*2]};
assign pixels_12_17 = {data_out[557*word_length*2-1 -: word_length*2]};
assign pixels_13_17 = {data_out[558*word_length*2-1 -: word_length*2]};
assign pixels_14_17 = {data_out[559*word_length*2-1 -: word_length*2]};
assign pixels_15_17 = {data_out[560*word_length*2-1 -: word_length*2]};
assign pixels_16_17 = {data_out[561*word_length*2-1 -: word_length*2]};
assign pixels_17_17 = {data_out[562*word_length*2-1 -: word_length*2]};
assign pixels_18_17 = {data_out[563*word_length*2-1 -: word_length*2]};
assign pixels_19_17 = {data_out[564*word_length*2-1 -: word_length*2]};
assign pixels_20_17 = {data_out[565*word_length*2-1 -: word_length*2]};
assign pixels_21_17 = {data_out[566*word_length*2-1 -: word_length*2]};
assign pixels_22_17 = {data_out[567*word_length*2-1 -: word_length*2]};
assign pixels_23_17 = {data_out[568*word_length*2-1 -: word_length*2]};
assign pixels_24_17 = {data_out[569*word_length*2-1 -: word_length*2]};
assign pixels_25_17 = {data_out[570*word_length*2-1 -: word_length*2]};
assign pixels_26_17 = {data_out[571*word_length*2-1 -: word_length*2]};
assign pixels_27_17 = {data_out[572*word_length*2-1 -: word_length*2]};
assign pixels_28_17 = {data_out[573*word_length*2-1 -: word_length*2]};
assign pixels_29_17 = {data_out[574*word_length*2-1 -: word_length*2]};
assign pixels_30_17 = {data_out[575*word_length*2-1 -: word_length*2]};
assign pixels_31_17 = {data_out[576*word_length*2-1 -: word_length*2]};
assign pixels_0_18 = {data_out[577*word_length*2-1 -: word_length*2]};
assign pixels_1_18 = {data_out[578*word_length*2-1 -: word_length*2]};
assign pixels_2_18 = {data_out[579*word_length*2-1 -: word_length*2]};
assign pixels_3_18 = {data_out[580*word_length*2-1 -: word_length*2]};
assign pixels_4_18 = {data_out[581*word_length*2-1 -: word_length*2]};
assign pixels_5_18 = {data_out[582*word_length*2-1 -: word_length*2]};
assign pixels_6_18 = {data_out[583*word_length*2-1 -: word_length*2]};
assign pixels_7_18 = {data_out[584*word_length*2-1 -: word_length*2]};
assign pixels_8_18 = {data_out[585*word_length*2-1 -: word_length*2]};
assign pixels_9_18 = {data_out[586*word_length*2-1 -: word_length*2]};
assign pixels_10_18 = {data_out[587*word_length*2-1 -: word_length*2]};
assign pixels_11_18 = {data_out[588*word_length*2-1 -: word_length*2]};
assign pixels_12_18 = {data_out[589*word_length*2-1 -: word_length*2]};
assign pixels_13_18 = {data_out[590*word_length*2-1 -: word_length*2]};
assign pixels_14_18 = {data_out[591*word_length*2-1 -: word_length*2]};
assign pixels_15_18 = {data_out[592*word_length*2-1 -: word_length*2]};
assign pixels_16_18 = {data_out[593*word_length*2-1 -: word_length*2]};
assign pixels_17_18 = {data_out[594*word_length*2-1 -: word_length*2]};
assign pixels_18_18 = {data_out[595*word_length*2-1 -: word_length*2]};
assign pixels_19_18 = {data_out[596*word_length*2-1 -: word_length*2]};
assign pixels_20_18 = {data_out[597*word_length*2-1 -: word_length*2]};
assign pixels_21_18 = {data_out[598*word_length*2-1 -: word_length*2]};
assign pixels_22_18 = {data_out[599*word_length*2-1 -: word_length*2]};
assign pixels_23_18 = {data_out[600*word_length*2-1 -: word_length*2]};
assign pixels_24_18 = {data_out[601*word_length*2-1 -: word_length*2]};
assign pixels_25_18 = {data_out[602*word_length*2-1 -: word_length*2]};
assign pixels_26_18 = {data_out[603*word_length*2-1 -: word_length*2]};
assign pixels_27_18 = {data_out[604*word_length*2-1 -: word_length*2]};
assign pixels_28_18 = {data_out[605*word_length*2-1 -: word_length*2]};
assign pixels_29_18 = {data_out[606*word_length*2-1 -: word_length*2]};
assign pixels_30_18 = {data_out[607*word_length*2-1 -: word_length*2]};
assign pixels_31_18 = {data_out[608*word_length*2-1 -: word_length*2]};
assign pixels_0_19 = {data_out[609*word_length*2-1 -: word_length*2]};
assign pixels_1_19 = {data_out[610*word_length*2-1 -: word_length*2]};
assign pixels_2_19 = {data_out[611*word_length*2-1 -: word_length*2]};
assign pixels_3_19 = {data_out[612*word_length*2-1 -: word_length*2]};
assign pixels_4_19 = {data_out[613*word_length*2-1 -: word_length*2]};
assign pixels_5_19 = {data_out[614*word_length*2-1 -: word_length*2]};
assign pixels_6_19 = {data_out[615*word_length*2-1 -: word_length*2]};
assign pixels_7_19 = {data_out[616*word_length*2-1 -: word_length*2]};
assign pixels_8_19 = {data_out[617*word_length*2-1 -: word_length*2]};
assign pixels_9_19 = {data_out[618*word_length*2-1 -: word_length*2]};
assign pixels_10_19 = {data_out[619*word_length*2-1 -: word_length*2]};
assign pixels_11_19 = {data_out[620*word_length*2-1 -: word_length*2]};
assign pixels_12_19 = {data_out[621*word_length*2-1 -: word_length*2]};
assign pixels_13_19 = {data_out[622*word_length*2-1 -: word_length*2]};
assign pixels_14_19 = {data_out[623*word_length*2-1 -: word_length*2]};
assign pixels_15_19 = {data_out[624*word_length*2-1 -: word_length*2]};
assign pixels_16_19 = {data_out[625*word_length*2-1 -: word_length*2]};
assign pixels_17_19 = {data_out[626*word_length*2-1 -: word_length*2]};
assign pixels_18_19 = {data_out[627*word_length*2-1 -: word_length*2]};
assign pixels_19_19 = {data_out[628*word_length*2-1 -: word_length*2]};
assign pixels_20_19 = {data_out[629*word_length*2-1 -: word_length*2]};
assign pixels_21_19 = {data_out[630*word_length*2-1 -: word_length*2]};
assign pixels_22_19 = {data_out[631*word_length*2-1 -: word_length*2]};
assign pixels_23_19 = {data_out[632*word_length*2-1 -: word_length*2]};
assign pixels_24_19 = {data_out[633*word_length*2-1 -: word_length*2]};
assign pixels_25_19 = {data_out[634*word_length*2-1 -: word_length*2]};
assign pixels_26_19 = {data_out[635*word_length*2-1 -: word_length*2]};
assign pixels_27_19 = {data_out[636*word_length*2-1 -: word_length*2]};
assign pixels_28_19 = {data_out[637*word_length*2-1 -: word_length*2]};
assign pixels_29_19 = {data_out[638*word_length*2-1 -: word_length*2]};
assign pixels_30_19 = {data_out[639*word_length*2-1 -: word_length*2]};
assign pixels_31_19 = {data_out[640*word_length*2-1 -: word_length*2]};
assign pixels_0_20 = {data_out[641*word_length*2-1 -: word_length*2]};
assign pixels_1_20 = {data_out[642*word_length*2-1 -: word_length*2]};
assign pixels_2_20 = {data_out[643*word_length*2-1 -: word_length*2]};
assign pixels_3_20 = {data_out[644*word_length*2-1 -: word_length*2]};
assign pixels_4_20 = {data_out[645*word_length*2-1 -: word_length*2]};
assign pixels_5_20 = {data_out[646*word_length*2-1 -: word_length*2]};
assign pixels_6_20 = {data_out[647*word_length*2-1 -: word_length*2]};
assign pixels_7_20 = {data_out[648*word_length*2-1 -: word_length*2]};
assign pixels_8_20 = {data_out[649*word_length*2-1 -: word_length*2]};
assign pixels_9_20 = {data_out[650*word_length*2-1 -: word_length*2]};
assign pixels_10_20 = {data_out[651*word_length*2-1 -: word_length*2]};
assign pixels_11_20 = {data_out[652*word_length*2-1 -: word_length*2]};
assign pixels_12_20 = {data_out[653*word_length*2-1 -: word_length*2]};
assign pixels_13_20 = {data_out[654*word_length*2-1 -: word_length*2]};
assign pixels_14_20 = {data_out[655*word_length*2-1 -: word_length*2]};
assign pixels_15_20 = {data_out[656*word_length*2-1 -: word_length*2]};
assign pixels_16_20 = {data_out[657*word_length*2-1 -: word_length*2]};
assign pixels_17_20 = {data_out[658*word_length*2-1 -: word_length*2]};
assign pixels_18_20 = {data_out[659*word_length*2-1 -: word_length*2]};
assign pixels_19_20 = {data_out[660*word_length*2-1 -: word_length*2]};
assign pixels_20_20 = {data_out[661*word_length*2-1 -: word_length*2]};
assign pixels_21_20 = {data_out[662*word_length*2-1 -: word_length*2]};
assign pixels_22_20 = {data_out[663*word_length*2-1 -: word_length*2]};
assign pixels_23_20 = {data_out[664*word_length*2-1 -: word_length*2]};
assign pixels_24_20 = {data_out[665*word_length*2-1 -: word_length*2]};
assign pixels_25_20 = {data_out[666*word_length*2-1 -: word_length*2]};
assign pixels_26_20 = {data_out[667*word_length*2-1 -: word_length*2]};
assign pixels_27_20 = {data_out[668*word_length*2-1 -: word_length*2]};
assign pixels_28_20 = {data_out[669*word_length*2-1 -: word_length*2]};
assign pixels_29_20 = {data_out[670*word_length*2-1 -: word_length*2]};
assign pixels_30_20 = {data_out[671*word_length*2-1 -: word_length*2]};
assign pixels_31_20 = {data_out[672*word_length*2-1 -: word_length*2]};
assign pixels_0_21 = {data_out[673*word_length*2-1 -: word_length*2]};
assign pixels_1_21 = {data_out[674*word_length*2-1 -: word_length*2]};
assign pixels_2_21 = {data_out[675*word_length*2-1 -: word_length*2]};
assign pixels_3_21 = {data_out[676*word_length*2-1 -: word_length*2]};
assign pixels_4_21 = {data_out[677*word_length*2-1 -: word_length*2]};
assign pixels_5_21 = {data_out[678*word_length*2-1 -: word_length*2]};
assign pixels_6_21 = {data_out[679*word_length*2-1 -: word_length*2]};
assign pixels_7_21 = {data_out[680*word_length*2-1 -: word_length*2]};
assign pixels_8_21 = {data_out[681*word_length*2-1 -: word_length*2]};
assign pixels_9_21 = {data_out[682*word_length*2-1 -: word_length*2]};
assign pixels_10_21 = {data_out[683*word_length*2-1 -: word_length*2]};
assign pixels_11_21 = {data_out[684*word_length*2-1 -: word_length*2]};
assign pixels_12_21 = {data_out[685*word_length*2-1 -: word_length*2]};
assign pixels_13_21 = {data_out[686*word_length*2-1 -: word_length*2]};
assign pixels_14_21 = {data_out[687*word_length*2-1 -: word_length*2]};
assign pixels_15_21 = {data_out[688*word_length*2-1 -: word_length*2]};
assign pixels_16_21 = {data_out[689*word_length*2-1 -: word_length*2]};
assign pixels_17_21 = {data_out[690*word_length*2-1 -: word_length*2]};
assign pixels_18_21 = {data_out[691*word_length*2-1 -: word_length*2]};
assign pixels_19_21 = {data_out[692*word_length*2-1 -: word_length*2]};
assign pixels_20_21 = {data_out[693*word_length*2-1 -: word_length*2]};
assign pixels_21_21 = {data_out[694*word_length*2-1 -: word_length*2]};
assign pixels_22_21 = {data_out[695*word_length*2-1 -: word_length*2]};
assign pixels_23_21 = {data_out[696*word_length*2-1 -: word_length*2]};
assign pixels_24_21 = {data_out[697*word_length*2-1 -: word_length*2]};
assign pixels_25_21 = {data_out[698*word_length*2-1 -: word_length*2]};
assign pixels_26_21 = {data_out[699*word_length*2-1 -: word_length*2]};
assign pixels_27_21 = {data_out[700*word_length*2-1 -: word_length*2]};
assign pixels_28_21 = {data_out[701*word_length*2-1 -: word_length*2]};
assign pixels_29_21 = {data_out[702*word_length*2-1 -: word_length*2]};
assign pixels_30_21 = {data_out[703*word_length*2-1 -: word_length*2]};
assign pixels_31_21 = {data_out[704*word_length*2-1 -: word_length*2]};
assign pixels_0_22 = {data_out[705*word_length*2-1 -: word_length*2]};
assign pixels_1_22 = {data_out[706*word_length*2-1 -: word_length*2]};
assign pixels_2_22 = {data_out[707*word_length*2-1 -: word_length*2]};
assign pixels_3_22 = {data_out[708*word_length*2-1 -: word_length*2]};
assign pixels_4_22 = {data_out[709*word_length*2-1 -: word_length*2]};
assign pixels_5_22 = {data_out[710*word_length*2-1 -: word_length*2]};
assign pixels_6_22 = {data_out[711*word_length*2-1 -: word_length*2]};
assign pixels_7_22 = {data_out[712*word_length*2-1 -: word_length*2]};
assign pixels_8_22 = {data_out[713*word_length*2-1 -: word_length*2]};
assign pixels_9_22 = {data_out[714*word_length*2-1 -: word_length*2]};
assign pixels_10_22 = {data_out[715*word_length*2-1 -: word_length*2]};
assign pixels_11_22 = {data_out[716*word_length*2-1 -: word_length*2]};
assign pixels_12_22 = {data_out[717*word_length*2-1 -: word_length*2]};
assign pixels_13_22 = {data_out[718*word_length*2-1 -: word_length*2]};
assign pixels_14_22 = {data_out[719*word_length*2-1 -: word_length*2]};
assign pixels_15_22 = {data_out[720*word_length*2-1 -: word_length*2]};
assign pixels_16_22 = {data_out[721*word_length*2-1 -: word_length*2]};
assign pixels_17_22 = {data_out[722*word_length*2-1 -: word_length*2]};
assign pixels_18_22 = {data_out[723*word_length*2-1 -: word_length*2]};
assign pixels_19_22 = {data_out[724*word_length*2-1 -: word_length*2]};
assign pixels_20_22 = {data_out[725*word_length*2-1 -: word_length*2]};
assign pixels_21_22 = {data_out[726*word_length*2-1 -: word_length*2]};
assign pixels_22_22 = {data_out[727*word_length*2-1 -: word_length*2]};
assign pixels_23_22 = {data_out[728*word_length*2-1 -: word_length*2]};
assign pixels_24_22 = {data_out[729*word_length*2-1 -: word_length*2]};
assign pixels_25_22 = {data_out[730*word_length*2-1 -: word_length*2]};
assign pixels_26_22 = {data_out[731*word_length*2-1 -: word_length*2]};
assign pixels_27_22 = {data_out[732*word_length*2-1 -: word_length*2]};
assign pixels_28_22 = {data_out[733*word_length*2-1 -: word_length*2]};
assign pixels_29_22 = {data_out[734*word_length*2-1 -: word_length*2]};
assign pixels_30_22 = {data_out[735*word_length*2-1 -: word_length*2]};
assign pixels_31_22 = {data_out[736*word_length*2-1 -: word_length*2]};
assign pixels_0_23 = {data_out[737*word_length*2-1 -: word_length*2]};
assign pixels_1_23 = {data_out[738*word_length*2-1 -: word_length*2]};
assign pixels_2_23 = {data_out[739*word_length*2-1 -: word_length*2]};
assign pixels_3_23 = {data_out[740*word_length*2-1 -: word_length*2]};
assign pixels_4_23 = {data_out[741*word_length*2-1 -: word_length*2]};
assign pixels_5_23 = {data_out[742*word_length*2-1 -: word_length*2]};
assign pixels_6_23 = {data_out[743*word_length*2-1 -: word_length*2]};
assign pixels_7_23 = {data_out[744*word_length*2-1 -: word_length*2]};
assign pixels_8_23 = {data_out[745*word_length*2-1 -: word_length*2]};
assign pixels_9_23 = {data_out[746*word_length*2-1 -: word_length*2]};
assign pixels_10_23 = {data_out[747*word_length*2-1 -: word_length*2]};
assign pixels_11_23 = {data_out[748*word_length*2-1 -: word_length*2]};
assign pixels_12_23 = {data_out[749*word_length*2-1 -: word_length*2]};
assign pixels_13_23 = {data_out[750*word_length*2-1 -: word_length*2]};
assign pixels_14_23 = {data_out[751*word_length*2-1 -: word_length*2]};
assign pixels_15_23 = {data_out[752*word_length*2-1 -: word_length*2]};
assign pixels_16_23 = {data_out[753*word_length*2-1 -: word_length*2]};
assign pixels_17_23 = {data_out[754*word_length*2-1 -: word_length*2]};
assign pixels_18_23 = {data_out[755*word_length*2-1 -: word_length*2]};
assign pixels_19_23 = {data_out[756*word_length*2-1 -: word_length*2]};
assign pixels_20_23 = {data_out[757*word_length*2-1 -: word_length*2]};
assign pixels_21_23 = {data_out[758*word_length*2-1 -: word_length*2]};
assign pixels_22_23 = {data_out[759*word_length*2-1 -: word_length*2]};
assign pixels_23_23 = {data_out[760*word_length*2-1 -: word_length*2]};
assign pixels_24_23 = {data_out[761*word_length*2-1 -: word_length*2]};
assign pixels_25_23 = {data_out[762*word_length*2-1 -: word_length*2]};
assign pixels_26_23 = {data_out[763*word_length*2-1 -: word_length*2]};
assign pixels_27_23 = {data_out[764*word_length*2-1 -: word_length*2]};
assign pixels_28_23 = {data_out[765*word_length*2-1 -: word_length*2]};
assign pixels_29_23 = {data_out[766*word_length*2-1 -: word_length*2]};
assign pixels_30_23 = {data_out[767*word_length*2-1 -: word_length*2]};
assign pixels_31_23 = {data_out[768*word_length*2-1 -: word_length*2]};
assign pixels_0_24 = {data_out[769*word_length*2-1 -: word_length*2]};
assign pixels_1_24 = {data_out[770*word_length*2-1 -: word_length*2]};
assign pixels_2_24 = {data_out[771*word_length*2-1 -: word_length*2]};
assign pixels_3_24 = {data_out[772*word_length*2-1 -: word_length*2]};
assign pixels_4_24 = {data_out[773*word_length*2-1 -: word_length*2]};
assign pixels_5_24 = {data_out[774*word_length*2-1 -: word_length*2]};
assign pixels_6_24 = {data_out[775*word_length*2-1 -: word_length*2]};
assign pixels_7_24 = {data_out[776*word_length*2-1 -: word_length*2]};
assign pixels_8_24 = {data_out[777*word_length*2-1 -: word_length*2]};
assign pixels_9_24 = {data_out[778*word_length*2-1 -: word_length*2]};
assign pixels_10_24 = {data_out[779*word_length*2-1 -: word_length*2]};
assign pixels_11_24 = {data_out[780*word_length*2-1 -: word_length*2]};
assign pixels_12_24 = {data_out[781*word_length*2-1 -: word_length*2]};
assign pixels_13_24 = {data_out[782*word_length*2-1 -: word_length*2]};
assign pixels_14_24 = {data_out[783*word_length*2-1 -: word_length*2]};
assign pixels_15_24 = {data_out[784*word_length*2-1 -: word_length*2]};
assign pixels_16_24 = {data_out[785*word_length*2-1 -: word_length*2]};
assign pixels_17_24 = {data_out[786*word_length*2-1 -: word_length*2]};
assign pixels_18_24 = {data_out[787*word_length*2-1 -: word_length*2]};
assign pixels_19_24 = {data_out[788*word_length*2-1 -: word_length*2]};
assign pixels_20_24 = {data_out[789*word_length*2-1 -: word_length*2]};
assign pixels_21_24 = {data_out[790*word_length*2-1 -: word_length*2]};
assign pixels_22_24 = {data_out[791*word_length*2-1 -: word_length*2]};
assign pixels_23_24 = {data_out[792*word_length*2-1 -: word_length*2]};
assign pixels_24_24 = {data_out[793*word_length*2-1 -: word_length*2]};
assign pixels_25_24 = {data_out[794*word_length*2-1 -: word_length*2]};
assign pixels_26_24 = {data_out[795*word_length*2-1 -: word_length*2]};
assign pixels_27_24 = {data_out[796*word_length*2-1 -: word_length*2]};
assign pixels_28_24 = {data_out[797*word_length*2-1 -: word_length*2]};
assign pixels_29_24 = {data_out[798*word_length*2-1 -: word_length*2]};
assign pixels_30_24 = {data_out[799*word_length*2-1 -: word_length*2]};
assign pixels_31_24 = {data_out[800*word_length*2-1 -: word_length*2]};
assign pixels_0_25 = {data_out[801*word_length*2-1 -: word_length*2]};
assign pixels_1_25 = {data_out[802*word_length*2-1 -: word_length*2]};
assign pixels_2_25 = {data_out[803*word_length*2-1 -: word_length*2]};
assign pixels_3_25 = {data_out[804*word_length*2-1 -: word_length*2]};
assign pixels_4_25 = {data_out[805*word_length*2-1 -: word_length*2]};
assign pixels_5_25 = {data_out[806*word_length*2-1 -: word_length*2]};
assign pixels_6_25 = {data_out[807*word_length*2-1 -: word_length*2]};
assign pixels_7_25 = {data_out[808*word_length*2-1 -: word_length*2]};
assign pixels_8_25 = {data_out[809*word_length*2-1 -: word_length*2]};
assign pixels_9_25 = {data_out[810*word_length*2-1 -: word_length*2]};
assign pixels_10_25 = {data_out[811*word_length*2-1 -: word_length*2]};
assign pixels_11_25 = {data_out[812*word_length*2-1 -: word_length*2]};
assign pixels_12_25 = {data_out[813*word_length*2-1 -: word_length*2]};
assign pixels_13_25 = {data_out[814*word_length*2-1 -: word_length*2]};
assign pixels_14_25 = {data_out[815*word_length*2-1 -: word_length*2]};
assign pixels_15_25 = {data_out[816*word_length*2-1 -: word_length*2]};
assign pixels_16_25 = {data_out[817*word_length*2-1 -: word_length*2]};
assign pixels_17_25 = {data_out[818*word_length*2-1 -: word_length*2]};
assign pixels_18_25 = {data_out[819*word_length*2-1 -: word_length*2]};
assign pixels_19_25 = {data_out[820*word_length*2-1 -: word_length*2]};
assign pixels_20_25 = {data_out[821*word_length*2-1 -: word_length*2]};
assign pixels_21_25 = {data_out[822*word_length*2-1 -: word_length*2]};
assign pixels_22_25 = {data_out[823*word_length*2-1 -: word_length*2]};
assign pixels_23_25 = {data_out[824*word_length*2-1 -: word_length*2]};
assign pixels_24_25 = {data_out[825*word_length*2-1 -: word_length*2]};
assign pixels_25_25 = {data_out[826*word_length*2-1 -: word_length*2]};
assign pixels_26_25 = {data_out[827*word_length*2-1 -: word_length*2]};
assign pixels_27_25 = {data_out[828*word_length*2-1 -: word_length*2]};
assign pixels_28_25 = {data_out[829*word_length*2-1 -: word_length*2]};
assign pixels_29_25 = {data_out[830*word_length*2-1 -: word_length*2]};
assign pixels_30_25 = {data_out[831*word_length*2-1 -: word_length*2]};
assign pixels_31_25 = {data_out[832*word_length*2-1 -: word_length*2]};
assign pixels_0_26 = {data_out[833*word_length*2-1 -: word_length*2]};
assign pixels_1_26 = {data_out[834*word_length*2-1 -: word_length*2]};
assign pixels_2_26 = {data_out[835*word_length*2-1 -: word_length*2]};
assign pixels_3_26 = {data_out[836*word_length*2-1 -: word_length*2]};
assign pixels_4_26 = {data_out[837*word_length*2-1 -: word_length*2]};
assign pixels_5_26 = {data_out[838*word_length*2-1 -: word_length*2]};
assign pixels_6_26 = {data_out[839*word_length*2-1 -: word_length*2]};
assign pixels_7_26 = {data_out[840*word_length*2-1 -: word_length*2]};
assign pixels_8_26 = {data_out[841*word_length*2-1 -: word_length*2]};
assign pixels_9_26 = {data_out[842*word_length*2-1 -: word_length*2]};
assign pixels_10_26 = {data_out[843*word_length*2-1 -: word_length*2]};
assign pixels_11_26 = {data_out[844*word_length*2-1 -: word_length*2]};
assign pixels_12_26 = {data_out[845*word_length*2-1 -: word_length*2]};
assign pixels_13_26 = {data_out[846*word_length*2-1 -: word_length*2]};
assign pixels_14_26 = {data_out[847*word_length*2-1 -: word_length*2]};
assign pixels_15_26 = {data_out[848*word_length*2-1 -: word_length*2]};
assign pixels_16_26 = {data_out[849*word_length*2-1 -: word_length*2]};
assign pixels_17_26 = {data_out[850*word_length*2-1 -: word_length*2]};
assign pixels_18_26 = {data_out[851*word_length*2-1 -: word_length*2]};
assign pixels_19_26 = {data_out[852*word_length*2-1 -: word_length*2]};
assign pixels_20_26 = {data_out[853*word_length*2-1 -: word_length*2]};
assign pixels_21_26 = {data_out[854*word_length*2-1 -: word_length*2]};
assign pixels_22_26 = {data_out[855*word_length*2-1 -: word_length*2]};
assign pixels_23_26 = {data_out[856*word_length*2-1 -: word_length*2]};
assign pixels_24_26 = {data_out[857*word_length*2-1 -: word_length*2]};
assign pixels_25_26 = {data_out[858*word_length*2-1 -: word_length*2]};
assign pixels_26_26 = {data_out[859*word_length*2-1 -: word_length*2]};
assign pixels_27_26 = {data_out[860*word_length*2-1 -: word_length*2]};
assign pixels_28_26 = {data_out[861*word_length*2-1 -: word_length*2]};
assign pixels_29_26 = {data_out[862*word_length*2-1 -: word_length*2]};
assign pixels_30_26 = {data_out[863*word_length*2-1 -: word_length*2]};
assign pixels_31_26 = {data_out[864*word_length*2-1 -: word_length*2]};
assign pixels_0_27 = {data_out[865*word_length*2-1 -: word_length*2]};
assign pixels_1_27 = {data_out[866*word_length*2-1 -: word_length*2]};
assign pixels_2_27 = {data_out[867*word_length*2-1 -: word_length*2]};
assign pixels_3_27 = {data_out[868*word_length*2-1 -: word_length*2]};
assign pixels_4_27 = {data_out[869*word_length*2-1 -: word_length*2]};
assign pixels_5_27 = {data_out[870*word_length*2-1 -: word_length*2]};
assign pixels_6_27 = {data_out[871*word_length*2-1 -: word_length*2]};
assign pixels_7_27 = {data_out[872*word_length*2-1 -: word_length*2]};
assign pixels_8_27 = {data_out[873*word_length*2-1 -: word_length*2]};
assign pixels_9_27 = {data_out[874*word_length*2-1 -: word_length*2]};
assign pixels_10_27 = {data_out[875*word_length*2-1 -: word_length*2]};
assign pixels_11_27 = {data_out[876*word_length*2-1 -: word_length*2]};
assign pixels_12_27 = {data_out[877*word_length*2-1 -: word_length*2]};
assign pixels_13_27 = {data_out[878*word_length*2-1 -: word_length*2]};
assign pixels_14_27 = {data_out[879*word_length*2-1 -: word_length*2]};
assign pixels_15_27 = {data_out[880*word_length*2-1 -: word_length*2]};
assign pixels_16_27 = {data_out[881*word_length*2-1 -: word_length*2]};
assign pixels_17_27 = {data_out[882*word_length*2-1 -: word_length*2]};
assign pixels_18_27 = {data_out[883*word_length*2-1 -: word_length*2]};
assign pixels_19_27 = {data_out[884*word_length*2-1 -: word_length*2]};
assign pixels_20_27 = {data_out[885*word_length*2-1 -: word_length*2]};
assign pixels_21_27 = {data_out[886*word_length*2-1 -: word_length*2]};
assign pixels_22_27 = {data_out[887*word_length*2-1 -: word_length*2]};
assign pixels_23_27 = {data_out[888*word_length*2-1 -: word_length*2]};
assign pixels_24_27 = {data_out[889*word_length*2-1 -: word_length*2]};
assign pixels_25_27 = {data_out[890*word_length*2-1 -: word_length*2]};
assign pixels_26_27 = {data_out[891*word_length*2-1 -: word_length*2]};
assign pixels_27_27 = {data_out[892*word_length*2-1 -: word_length*2]};
assign pixels_28_27 = {data_out[893*word_length*2-1 -: word_length*2]};
assign pixels_29_27 = {data_out[894*word_length*2-1 -: word_length*2]};
assign pixels_30_27 = {data_out[895*word_length*2-1 -: word_length*2]};
assign pixels_31_27 = {data_out[896*word_length*2-1 -: word_length*2]};
assign pixels_0_28 = {data_out[897*word_length*2-1 -: word_length*2]};
assign pixels_1_28 = {data_out[898*word_length*2-1 -: word_length*2]};
assign pixels_2_28 = {data_out[899*word_length*2-1 -: word_length*2]};
assign pixels_3_28 = {data_out[900*word_length*2-1 -: word_length*2]};
assign pixels_4_28 = {data_out[901*word_length*2-1 -: word_length*2]};
assign pixels_5_28 = {data_out[902*word_length*2-1 -: word_length*2]};
assign pixels_6_28 = {data_out[903*word_length*2-1 -: word_length*2]};
assign pixels_7_28 = {data_out[904*word_length*2-1 -: word_length*2]};
assign pixels_8_28 = {data_out[905*word_length*2-1 -: word_length*2]};
assign pixels_9_28 = {data_out[906*word_length*2-1 -: word_length*2]};
assign pixels_10_28 = {data_out[907*word_length*2-1 -: word_length*2]};
assign pixels_11_28 = {data_out[908*word_length*2-1 -: word_length*2]};
assign pixels_12_28 = {data_out[909*word_length*2-1 -: word_length*2]};
assign pixels_13_28 = {data_out[910*word_length*2-1 -: word_length*2]};
assign pixels_14_28 = {data_out[911*word_length*2-1 -: word_length*2]};
assign pixels_15_28 = {data_out[912*word_length*2-1 -: word_length*2]};
assign pixels_16_28 = {data_out[913*word_length*2-1 -: word_length*2]};
assign pixels_17_28 = {data_out[914*word_length*2-1 -: word_length*2]};
assign pixels_18_28 = {data_out[915*word_length*2-1 -: word_length*2]};
assign pixels_19_28 = {data_out[916*word_length*2-1 -: word_length*2]};
assign pixels_20_28 = {data_out[917*word_length*2-1 -: word_length*2]};
assign pixels_21_28 = {data_out[918*word_length*2-1 -: word_length*2]};
assign pixels_22_28 = {data_out[919*word_length*2-1 -: word_length*2]};
assign pixels_23_28 = {data_out[920*word_length*2-1 -: word_length*2]};
assign pixels_24_28 = {data_out[921*word_length*2-1 -: word_length*2]};
assign pixels_25_28 = {data_out[922*word_length*2-1 -: word_length*2]};
assign pixels_26_28 = {data_out[923*word_length*2-1 -: word_length*2]};
assign pixels_27_28 = {data_out[924*word_length*2-1 -: word_length*2]};
assign pixels_28_28 = {data_out[925*word_length*2-1 -: word_length*2]};
assign pixels_29_28 = {data_out[926*word_length*2-1 -: word_length*2]};
assign pixels_30_28 = {data_out[927*word_length*2-1 -: word_length*2]};
assign pixels_31_28 = {data_out[928*word_length*2-1 -: word_length*2]};
assign pixels_0_29 = {data_out[929*word_length*2-1 -: word_length*2]};
assign pixels_1_29 = {data_out[930*word_length*2-1 -: word_length*2]};
assign pixels_2_29 = {data_out[931*word_length*2-1 -: word_length*2]};
assign pixels_3_29 = {data_out[932*word_length*2-1 -: word_length*2]};
assign pixels_4_29 = {data_out[933*word_length*2-1 -: word_length*2]};
assign pixels_5_29 = {data_out[934*word_length*2-1 -: word_length*2]};
assign pixels_6_29 = {data_out[935*word_length*2-1 -: word_length*2]};
assign pixels_7_29 = {data_out[936*word_length*2-1 -: word_length*2]};
assign pixels_8_29 = {data_out[937*word_length*2-1 -: word_length*2]};
assign pixels_9_29 = {data_out[938*word_length*2-1 -: word_length*2]};
assign pixels_10_29 = {data_out[939*word_length*2-1 -: word_length*2]};
assign pixels_11_29 = {data_out[940*word_length*2-1 -: word_length*2]};
assign pixels_12_29 = {data_out[941*word_length*2-1 -: word_length*2]};
assign pixels_13_29 = {data_out[942*word_length*2-1 -: word_length*2]};
assign pixels_14_29 = {data_out[943*word_length*2-1 -: word_length*2]};
assign pixels_15_29 = {data_out[944*word_length*2-1 -: word_length*2]};
assign pixels_16_29 = {data_out[945*word_length*2-1 -: word_length*2]};
assign pixels_17_29 = {data_out[946*word_length*2-1 -: word_length*2]};
assign pixels_18_29 = {data_out[947*word_length*2-1 -: word_length*2]};
assign pixels_19_29 = {data_out[948*word_length*2-1 -: word_length*2]};
assign pixels_20_29 = {data_out[949*word_length*2-1 -: word_length*2]};
assign pixels_21_29 = {data_out[950*word_length*2-1 -: word_length*2]};
assign pixels_22_29 = {data_out[951*word_length*2-1 -: word_length*2]};
assign pixels_23_29 = {data_out[952*word_length*2-1 -: word_length*2]};
assign pixels_24_29 = {data_out[953*word_length*2-1 -: word_length*2]};
assign pixels_25_29 = {data_out[954*word_length*2-1 -: word_length*2]};
assign pixels_26_29 = {data_out[955*word_length*2-1 -: word_length*2]};
assign pixels_27_29 = {data_out[956*word_length*2-1 -: word_length*2]};
assign pixels_28_29 = {data_out[957*word_length*2-1 -: word_length*2]};
assign pixels_29_29 = {data_out[958*word_length*2-1 -: word_length*2]};
assign pixels_30_29 = {data_out[959*word_length*2-1 -: word_length*2]};
assign pixels_31_29 = {data_out[960*word_length*2-1 -: word_length*2]};
assign pixels_0_30 = {data_out[961*word_length*2-1 -: word_length*2]};
assign pixels_1_30 = {data_out[962*word_length*2-1 -: word_length*2]};
assign pixels_2_30 = {data_out[963*word_length*2-1 -: word_length*2]};
assign pixels_3_30 = {data_out[964*word_length*2-1 -: word_length*2]};
assign pixels_4_30 = {data_out[965*word_length*2-1 -: word_length*2]};
assign pixels_5_30 = {data_out[966*word_length*2-1 -: word_length*2]};
assign pixels_6_30 = {data_out[967*word_length*2-1 -: word_length*2]};
assign pixels_7_30 = {data_out[968*word_length*2-1 -: word_length*2]};
assign pixels_8_30 = {data_out[969*word_length*2-1 -: word_length*2]};
assign pixels_9_30 = {data_out[970*word_length*2-1 -: word_length*2]};
assign pixels_10_30 = {data_out[971*word_length*2-1 -: word_length*2]};
assign pixels_11_30 = {data_out[972*word_length*2-1 -: word_length*2]};
assign pixels_12_30 = {data_out[973*word_length*2-1 -: word_length*2]};
assign pixels_13_30 = {data_out[974*word_length*2-1 -: word_length*2]};
assign pixels_14_30 = {data_out[975*word_length*2-1 -: word_length*2]};
assign pixels_15_30 = {data_out[976*word_length*2-1 -: word_length*2]};
assign pixels_16_30 = {data_out[977*word_length*2-1 -: word_length*2]};
assign pixels_17_30 = {data_out[978*word_length*2-1 -: word_length*2]};
assign pixels_18_30 = {data_out[979*word_length*2-1 -: word_length*2]};
assign pixels_19_30 = {data_out[980*word_length*2-1 -: word_length*2]};
assign pixels_20_30 = {data_out[981*word_length*2-1 -: word_length*2]};
assign pixels_21_30 = {data_out[982*word_length*2-1 -: word_length*2]};
assign pixels_22_30 = {data_out[983*word_length*2-1 -: word_length*2]};
assign pixels_23_30 = {data_out[984*word_length*2-1 -: word_length*2]};
assign pixels_24_30 = {data_out[985*word_length*2-1 -: word_length*2]};
assign pixels_25_30 = {data_out[986*word_length*2-1 -: word_length*2]};
assign pixels_26_30 = {data_out[987*word_length*2-1 -: word_length*2]};
assign pixels_27_30 = {data_out[988*word_length*2-1 -: word_length*2]};
assign pixels_28_30 = {data_out[989*word_length*2-1 -: word_length*2]};
assign pixels_29_30 = {data_out[990*word_length*2-1 -: word_length*2]};
assign pixels_30_30 = {data_out[991*word_length*2-1 -: word_length*2]};
assign pixels_31_30 = {data_out[992*word_length*2-1 -: word_length*2]};
assign pixels_0_31 = {data_out[993*word_length*2-1 -: word_length*2]};
assign pixels_1_31 = {data_out[994*word_length*2-1 -: word_length*2]};
assign pixels_2_31 = {data_out[995*word_length*2-1 -: word_length*2]};
assign pixels_3_31 = {data_out[996*word_length*2-1 -: word_length*2]};
assign pixels_4_31 = {data_out[997*word_length*2-1 -: word_length*2]};
assign pixels_5_31 = {data_out[998*word_length*2-1 -: word_length*2]};
assign pixels_6_31 = {data_out[999*word_length*2-1 -: word_length*2]};
assign pixels_7_31 = {data_out[1000*word_length*2-1 -: word_length*2]};
assign pixels_8_31 = {data_out[1001*word_length*2-1 -: word_length*2]};
assign pixels_9_31 = {data_out[1002*word_length*2-1 -: word_length*2]};
assign pixels_10_31 = {data_out[1003*word_length*2-1 -: word_length*2]};
assign pixels_11_31 = {data_out[1004*word_length*2-1 -: word_length*2]};
assign pixels_12_31 = {data_out[1005*word_length*2-1 -: word_length*2]};
assign pixels_13_31 = {data_out[1006*word_length*2-1 -: word_length*2]};
assign pixels_14_31 = {data_out[1007*word_length*2-1 -: word_length*2]};
assign pixels_15_31 = {data_out[1008*word_length*2-1 -: word_length*2]};
assign pixels_16_31 = {data_out[1009*word_length*2-1 -: word_length*2]};
assign pixels_17_31 = {data_out[1010*word_length*2-1 -: word_length*2]};
assign pixels_18_31 = {data_out[1011*word_length*2-1 -: word_length*2]};
assign pixels_19_31 = {data_out[1012*word_length*2-1 -: word_length*2]};
assign pixels_20_31 = {data_out[1013*word_length*2-1 -: word_length*2]};
assign pixels_21_31 = {data_out[1014*word_length*2-1 -: word_length*2]};
assign pixels_22_31 = {data_out[1015*word_length*2-1 -: word_length*2]};
assign pixels_23_31 = {data_out[1016*word_length*2-1 -: word_length*2]};
assign pixels_24_31 = {data_out[1017*word_length*2-1 -: word_length*2]};
assign pixels_25_31 = {data_out[1018*word_length*2-1 -: word_length*2]};
assign pixels_26_31 = {data_out[1019*word_length*2-1 -: word_length*2]};
assign pixels_27_31 = {data_out[1020*word_length*2-1 -: word_length*2]};
assign pixels_28_31 = {data_out[1021*word_length*2-1 -: word_length*2]};
assign pixels_29_31 = {data_out[1022*word_length*2-1 -: word_length*2]};
assign pixels_30_31 = {data_out[1023*word_length*2-1 -: word_length*2]};
assign pixels_31_31 = {data_out[1024*word_length*2-1 -: word_length*2]};


//iter
integer i;

initial begin
    #0      rst = 0;
            clk = 1;
            weight_value = 'h19_05_00_0b_fc_ed_12_f6_02_f7_08_0d_05_dd_fc_ed_f1_ff_09_fa_00_07_f2_ee_e7;
            //weight_value = {25{16'h0010}};
    #10     rst = 1;
    #10     rst = 0;
    #100    in_valid = 1;
            for (i=0;i<(image_size*image_size);i=i+1)begin
                data_in[word_length-1:0] = {pe_input_feature_value[(i+1)*word_length-1 -:word_length]};
                //data_in[word_length-1:0] = i+1;
                #10;
            end
    #1000;
    if(pixels_0_0!==16'hff1f) $display("ERROR! at (0,0)\n");
if(pixels_1_0!==16'h0195) $display("ERROR! at (1,0)\n");
if(pixels_2_0!==16'hfe66) $display("ERROR! at (2,0)\n");
if(pixels_3_0!==16'hffe8) $display("ERROR! at (3,0)\n");
if(pixels_4_0!==16'h00db) $display("ERROR! at (4,0)\n");
if(pixels_5_0!==16'hff04) $display("ERROR! at (5,0)\n");
if(pixels_6_0!==16'h013d) $display("ERROR! at (6,0)\n");
if(pixels_7_0!==16'hfec0) $display("ERROR! at (7,0)\n");
if(pixels_8_0!==16'h02e9) $display("ERROR! at (8,0)\n");
if(pixels_9_0!==16'h008a) $display("ERROR! at (9,0)\n");
if(pixels_10_0!==16'h009a) $display("ERROR! at (10,0)\n");
if(pixels_11_0!==16'h049b) $display("ERROR! at (11,0)\n");
if(pixels_12_0!==16'hfff4) $display("ERROR! at (12,0)\n");
if(pixels_13_0!==16'h009b) $display("ERROR! at (13,0)\n");
if(pixels_14_0!==16'hff7b) $display("ERROR! at (14,0)\n");
if(pixels_15_0!==16'hff55) $display("ERROR! at (15,0)\n");
if(pixels_16_0!==16'h009b) $display("ERROR! at (16,0)\n");
if(pixels_17_0!==16'h02c0) $display("ERROR! at (17,0)\n");
if(pixels_18_0!==16'h01ef) $display("ERROR! at (18,0)\n");
if(pixels_19_0!==16'hff44) $display("ERROR! at (19,0)\n");
if(pixels_20_0!==16'hfff6) $display("ERROR! at (20,0)\n");
if(pixels_21_0!==16'h000e) $display("ERROR! at (21,0)\n");
if(pixels_22_0!==16'hfc61) $display("ERROR! at (22,0)\n");
if(pixels_23_0!==16'h01ff) $display("ERROR! at (23,0)\n");
if(pixels_24_0!==16'hffc6) $display("ERROR! at (24,0)\n");
if(pixels_25_0!==16'hff8b) $display("ERROR! at (25,0)\n");
if(pixels_26_0!==16'h0761) $display("ERROR! at (26,0)\n");
if(pixels_27_0!==16'h0049) $display("ERROR! at (27,0)\n");
if(pixels_28_0!==16'h00be) $display("ERROR! at (28,0)\n");
if(pixels_29_0!==16'h022d) $display("ERROR! at (29,0)\n");
if(pixels_30_0!==16'hff3a) $display("ERROR! at (30,0)\n");
if(pixels_31_0!==16'hfff8) $display("ERROR! at (31,0)\n");
if(pixels_0_1!==16'h0209) $display("ERROR! at (0,1)\n");
if(pixels_1_1!==16'hfcbe) $display("ERROR! at (1,1)\n");
if(pixels_2_1!==16'h0266) $display("ERROR! at (2,1)\n");
if(pixels_3_1!==16'hfc11) $display("ERROR! at (3,1)\n");
if(pixels_4_1!==16'h0022) $display("ERROR! at (4,1)\n");
if(pixels_5_1!==16'hfe3d) $display("ERROR! at (5,1)\n");
if(pixels_6_1!==16'h0536) $display("ERROR! at (6,1)\n");
if(pixels_7_1!==16'h0079) $display("ERROR! at (7,1)\n");
if(pixels_8_1!==16'hfa9f) $display("ERROR! at (8,1)\n");
if(pixels_9_1!==16'h0579) $display("ERROR! at (9,1)\n");
if(pixels_10_1!==16'hfb9b) $display("ERROR! at (10,1)\n");
if(pixels_11_1!==16'h0081) $display("ERROR! at (11,1)\n");
if(pixels_12_1!==16'h01e0) $display("ERROR! at (12,1)\n");
if(pixels_13_1!==16'hfef3) $display("ERROR! at (13,1)\n");
if(pixels_14_1!==16'h0472) $display("ERROR! at (14,1)\n");
if(pixels_15_1!==16'hfd25) $display("ERROR! at (15,1)\n");
if(pixels_16_1!==16'hfff1) $display("ERROR! at (16,1)\n");
if(pixels_17_1!==16'hff1d) $display("ERROR! at (17,1)\n");
if(pixels_18_1!==16'h03a1) $display("ERROR! at (18,1)\n");
if(pixels_19_1!==16'h0126) $display("ERROR! at (19,1)\n");
if(pixels_20_1!==16'hff77) $display("ERROR! at (20,1)\n");
if(pixels_21_1!==16'hff1a) $display("ERROR! at (21,1)\n");
if(pixels_22_1!==16'h0488) $display("ERROR! at (22,1)\n");
if(pixels_23_1!==16'hfb9a) $display("ERROR! at (23,1)\n");
if(pixels_24_1!==16'h02ac) $display("ERROR! at (24,1)\n");
if(pixels_25_1!==16'h000a) $display("ERROR! at (25,1)\n");
if(pixels_26_1!==16'h0040) $display("ERROR! at (26,1)\n");
if(pixels_27_1!==16'h0040) $display("ERROR! at (27,1)\n");
if(pixels_28_1!==16'hffac) $display("ERROR! at (28,1)\n");
if(pixels_29_1!==16'h0048) $display("ERROR! at (29,1)\n");
if(pixels_30_1!==16'hfd28) $display("ERROR! at (30,1)\n");
if(pixels_31_1!==16'h002a) $display("ERROR! at (31,1)\n");
if(pixels_0_2!==16'hfbc0) $display("ERROR! at (0,2)\n");
if(pixels_1_2!==16'hfedc) $display("ERROR! at (1,2)\n");
if(pixels_2_2!==16'hfcce) $display("ERROR! at (2,2)\n");
if(pixels_3_2!==16'h0009) $display("ERROR! at (3,2)\n");
if(pixels_4_2!==16'hfc86) $display("ERROR! at (4,2)\n");
if(pixels_5_2!==16'h038b) $display("ERROR! at (5,2)\n");
if(pixels_6_2!==16'hfae6) $display("ERROR! at (6,2)\n");
if(pixels_7_2!==16'h07a3) $display("ERROR! at (7,2)\n");
if(pixels_8_2!==16'hfe7e) $display("ERROR! at (8,2)\n");
if(pixels_9_2!==16'h01ac) $display("ERROR! at (9,2)\n");
if(pixels_10_2!==16'h0314) $display("ERROR! at (10,2)\n");
if(pixels_11_2!==16'hfc95) $display("ERROR! at (11,2)\n");
if(pixels_12_2!==16'h05a8) $display("ERROR! at (12,2)\n");
if(pixels_13_2!==16'h03c8) $display("ERROR! at (13,2)\n");
if(pixels_14_2!==16'hf92c) $display("ERROR! at (14,2)\n");
if(pixels_15_2!==16'h046d) $display("ERROR! at (15,2)\n");
if(pixels_16_2!==16'hff17) $display("ERROR! at (16,2)\n");
if(pixels_17_2!==16'h0386) $display("ERROR! at (17,2)\n");
if(pixels_18_2!==16'h0132) $display("ERROR! at (18,2)\n");
if(pixels_19_2!==16'h00b2) $display("ERROR! at (19,2)\n");
if(pixels_20_2!==16'hf965) $display("ERROR! at (20,2)\n");
if(pixels_21_2!==16'hfb33) $display("ERROR! at (21,2)\n");
if(pixels_22_2!==16'hfd7f) $display("ERROR! at (22,2)\n");
if(pixels_23_2!==16'h0201) $display("ERROR! at (23,2)\n");
if(pixels_24_2!==16'hfbca) $display("ERROR! at (24,2)\n");
if(pixels_25_2!==16'h0134) $display("ERROR! at (25,2)\n");
if(pixels_26_2!==16'hff39) $display("ERROR! at (26,2)\n");
if(pixels_27_2!==16'h068e) $display("ERROR! at (27,2)\n");
if(pixels_28_2!==16'hff79) $display("ERROR! at (28,2)\n");
if(pixels_29_2!==16'hf8c3) $display("ERROR! at (29,2)\n");
if(pixels_30_2!==16'hfebb) $display("ERROR! at (30,2)\n");
if(pixels_31_2!==16'h0033) $display("ERROR! at (31,2)\n");
if(pixels_0_3!==16'h030a) $display("ERROR! at (0,3)\n");
if(pixels_1_3!==16'h0189) $display("ERROR! at (1,3)\n");
if(pixels_2_3!==16'hffea) $display("ERROR! at (2,3)\n");
if(pixels_3_3!==16'hfbd9) $display("ERROR! at (3,3)\n");
if(pixels_4_3!==16'h0297) $display("ERROR! at (4,3)\n");
if(pixels_5_3!==16'hff42) $display("ERROR! at (5,3)\n");
if(pixels_6_3!==16'h0077) $display("ERROR! at (6,3)\n");
if(pixels_7_3!==16'h02ba) $display("ERROR! at (7,3)\n");
if(pixels_8_3!==16'hff85) $display("ERROR! at (8,3)\n");
if(pixels_9_3!==16'hf4f2) $display("ERROR! at (9,3)\n");
if(pixels_10_3!==16'hff05) $display("ERROR! at (10,3)\n");
if(pixels_11_3!==16'h03f6) $display("ERROR! at (11,3)\n");
if(pixels_12_3!==16'hfcf1) $display("ERROR! at (12,3)\n");
if(pixels_13_3!==16'hfd41) $display("ERROR! at (13,3)\n");
if(pixels_14_3!==16'h0223) $display("ERROR! at (14,3)\n");
if(pixels_15_3!==16'hfbce) $display("ERROR! at (15,3)\n");
if(pixels_16_3!==16'h039c) $display("ERROR! at (16,3)\n");
if(pixels_17_3!==16'hf3ef) $display("ERROR! at (17,3)\n");
if(pixels_18_3!==16'hfe5e) $display("ERROR! at (18,3)\n");
if(pixels_19_3!==16'h022e) $display("ERROR! at (19,3)\n");
if(pixels_20_3!==16'h0294) $display("ERROR! at (20,3)\n");
if(pixels_21_3!==16'hfb7d) $display("ERROR! at (21,3)\n");
if(pixels_22_3!==16'h013b) $display("ERROR! at (22,3)\n");
if(pixels_23_3!==16'h050b) $display("ERROR! at (23,3)\n");
if(pixels_24_3!==16'h000b) $display("ERROR! at (24,3)\n");
if(pixels_25_3!==16'hfbec) $display("ERROR! at (25,3)\n");
if(pixels_26_3!==16'hfb98) $display("ERROR! at (26,3)\n");
if(pixels_27_3!==16'h01f1) $display("ERROR! at (27,3)\n");
if(pixels_28_3!==16'hfe92) $display("ERROR! at (28,3)\n");
if(pixels_29_3!==16'hfd4e) $display("ERROR! at (29,3)\n");
if(pixels_30_3!==16'h01c2) $display("ERROR! at (30,3)\n");
if(pixels_31_3!==16'hff15) $display("ERROR! at (31,3)\n");
if(pixels_0_4!==16'hfea3) $display("ERROR! at (0,4)\n");
if(pixels_1_4!==16'hfbd4) $display("ERROR! at (1,4)\n");
if(pixels_2_4!==16'h0100) $display("ERROR! at (2,4)\n");
if(pixels_3_4!==16'h0489) $display("ERROR! at (3,4)\n");
if(pixels_4_4!==16'h053c) $display("ERROR! at (4,4)\n");
if(pixels_5_4!==16'h040f) $display("ERROR! at (5,4)\n");
if(pixels_6_4!==16'h027b) $display("ERROR! at (6,4)\n");
if(pixels_7_4!==16'hfe06) $display("ERROR! at (7,4)\n");
if(pixels_8_4!==16'h00cf) $display("ERROR! at (8,4)\n");
if(pixels_9_4!==16'h0814) $display("ERROR! at (9,4)\n");
if(pixels_10_4!==16'hfb6a) $display("ERROR! at (10,4)\n");
if(pixels_11_4!==16'hf9b6) $display("ERROR! at (11,4)\n");
if(pixels_12_4!==16'hfe46) $display("ERROR! at (12,4)\n");
if(pixels_13_4!==16'hfda1) $display("ERROR! at (13,4)\n");
if(pixels_14_4!==16'hfddf) $display("ERROR! at (14,4)\n");
if(pixels_15_4!==16'hfa96) $display("ERROR! at (15,4)\n");
if(pixels_16_4!==16'hfa06) $display("ERROR! at (16,4)\n");
if(pixels_17_4!==16'h079b) $display("ERROR! at (17,4)\n");
if(pixels_18_4!==16'hfe66) $display("ERROR! at (18,4)\n");
if(pixels_19_4!==16'hfe56) $display("ERROR! at (19,4)\n");
if(pixels_20_4!==16'hfb4c) $display("ERROR! at (20,4)\n");
if(pixels_21_4!==16'h000c) $display("ERROR! at (21,4)\n");
if(pixels_22_4!==16'hfd82) $display("ERROR! at (22,4)\n");
if(pixels_23_4!==16'h0395) $display("ERROR! at (23,4)\n");
if(pixels_24_4!==16'h079e) $display("ERROR! at (24,4)\n");
if(pixels_25_4!==16'h015d) $display("ERROR! at (25,4)\n");
if(pixels_26_4!==16'hfdcb) $display("ERROR! at (26,4)\n");
if(pixels_27_4!==16'h01d7) $display("ERROR! at (27,4)\n");
if(pixels_28_4!==16'h0430) $display("ERROR! at (28,4)\n");
if(pixels_29_4!==16'hf822) $display("ERROR! at (29,4)\n");
if(pixels_30_4!==16'hf78b) $display("ERROR! at (30,4)\n");
if(pixels_31_4!==16'hfef8) $display("ERROR! at (31,4)\n");
if(pixels_0_5!==16'h00dc) $display("ERROR! at (0,5)\n");
if(pixels_1_5!==16'h05ac) $display("ERROR! at (1,5)\n");
if(pixels_2_5!==16'h024d) $display("ERROR! at (2,5)\n");
if(pixels_3_5!==16'h0103) $display("ERROR! at (3,5)\n");
if(pixels_4_5!==16'hfcc4) $display("ERROR! at (4,5)\n");
if(pixels_5_5!==16'h042e) $display("ERROR! at (5,5)\n");
if(pixels_6_5!==16'h02a7) $display("ERROR! at (6,5)\n");
if(pixels_7_5!==16'h0301) $display("ERROR! at (7,5)\n");
if(pixels_8_5!==16'h005c) $display("ERROR! at (8,5)\n");
if(pixels_9_5!==16'h0191) $display("ERROR! at (9,5)\n");
if(pixels_10_5!==16'hfeed) $display("ERROR! at (10,5)\n");
if(pixels_11_5!==16'h000e) $display("ERROR! at (11,5)\n");
if(pixels_12_5!==16'hfac6) $display("ERROR! at (12,5)\n");
if(pixels_13_5!==16'h02e3) $display("ERROR! at (13,5)\n");
if(pixels_14_5!==16'hfaa9) $display("ERROR! at (14,5)\n");
if(pixels_15_5!==16'hf877) $display("ERROR! at (15,5)\n");
if(pixels_16_5!==16'h05b4) $display("ERROR! at (16,5)\n");
if(pixels_17_5!==16'h008c) $display("ERROR! at (17,5)\n");
if(pixels_18_5!==16'hfea0) $display("ERROR! at (18,5)\n");
if(pixels_19_5!==16'hfdd9) $display("ERROR! at (19,5)\n");
if(pixels_20_5!==16'h0053) $display("ERROR! at (20,5)\n");
if(pixels_21_5!==16'hffd0) $display("ERROR! at (21,5)\n");
if(pixels_22_5!==16'hfeb5) $display("ERROR! at (22,5)\n");
if(pixels_23_5!==16'h020d) $display("ERROR! at (23,5)\n");
if(pixels_24_5!==16'h0410) $display("ERROR! at (24,5)\n");
if(pixels_25_5!==16'h01f8) $display("ERROR! at (25,5)\n");
if(pixels_26_5!==16'hfbe6) $display("ERROR! at (26,5)\n");
if(pixels_27_5!==16'hffcc) $display("ERROR! at (27,5)\n");
if(pixels_28_5!==16'hff58) $display("ERROR! at (28,5)\n");
if(pixels_29_5!==16'h0012) $display("ERROR! at (29,5)\n");
if(pixels_30_5!==16'hfd63) $display("ERROR! at (30,5)\n");
if(pixels_31_5!==16'h007f) $display("ERROR! at (31,5)\n");
if(pixels_0_6!==16'h01df) $display("ERROR! at (0,6)\n");
if(pixels_1_6!==16'hfc3e) $display("ERROR! at (1,6)\n");
if(pixels_2_6!==16'h0041) $display("ERROR! at (2,6)\n");
if(pixels_3_6!==16'h00ff) $display("ERROR! at (3,6)\n");
if(pixels_4_6!==16'h05d3) $display("ERROR! at (4,6)\n");
if(pixels_5_6!==16'h0749) $display("ERROR! at (5,6)\n");
if(pixels_6_6!==16'h0323) $display("ERROR! at (6,6)\n");
if(pixels_7_6!==16'h0238) $display("ERROR! at (7,6)\n");
if(pixels_8_6!==16'h0138) $display("ERROR! at (8,6)\n");
if(pixels_9_6!==16'hfc89) $display("ERROR! at (9,6)\n");
if(pixels_10_6!==16'hfea3) $display("ERROR! at (10,6)\n");
if(pixels_11_6!==16'h0239) $display("ERROR! at (11,6)\n");
if(pixels_12_6!==16'hfa66) $display("ERROR! at (12,6)\n");
if(pixels_13_6!==16'hfc29) $display("ERROR! at (13,6)\n");
if(pixels_14_6!==16'h0a32) $display("ERROR! at (14,6)\n");
if(pixels_15_6!==16'hf7df) $display("ERROR! at (15,6)\n");
if(pixels_16_6!==16'hf45c) $display("ERROR! at (16,6)\n");
if(pixels_17_6!==16'hfe01) $display("ERROR! at (17,6)\n");
if(pixels_18_6!==16'hfe2e) $display("ERROR! at (18,6)\n");
if(pixels_19_6!==16'h0537) $display("ERROR! at (19,6)\n");
if(pixels_20_6!==16'hfadd) $display("ERROR! at (20,6)\n");
if(pixels_21_6!==16'h041b) $display("ERROR! at (21,6)\n");
if(pixels_22_6!==16'hfe78) $display("ERROR! at (22,6)\n");
if(pixels_23_6!==16'h02bb) $display("ERROR! at (23,6)\n");
if(pixels_24_6!==16'hfb89) $display("ERROR! at (24,6)\n");
if(pixels_25_6!==16'h03fa) $display("ERROR! at (25,6)\n");
if(pixels_26_6!==16'h0697) $display("ERROR! at (26,6)\n");
if(pixels_27_6!==16'hfe32) $display("ERROR! at (27,6)\n");
if(pixels_28_6!==16'h011e) $display("ERROR! at (28,6)\n");
if(pixels_29_6!==16'hfdbf) $display("ERROR! at (29,6)\n");
if(pixels_30_6!==16'h00d0) $display("ERROR! at (30,6)\n");
if(pixels_31_6!==16'hfcae) $display("ERROR! at (31,6)\n");
if(pixels_0_7!==16'hfeb3) $display("ERROR! at (0,7)\n");
if(pixels_1_7!==16'hfee5) $display("ERROR! at (1,7)\n");
if(pixels_2_7!==16'h02c5) $display("ERROR! at (2,7)\n");
if(pixels_3_7!==16'h0238) $display("ERROR! at (3,7)\n");
if(pixels_4_7!==16'hff23) $display("ERROR! at (4,7)\n");
if(pixels_5_7!==16'hfd4a) $display("ERROR! at (5,7)\n");
if(pixels_6_7!==16'h0537) $display("ERROR! at (6,7)\n");
if(pixels_7_7!==16'hf94b) $display("ERROR! at (7,7)\n");
if(pixels_8_7!==16'hfca3) $display("ERROR! at (8,7)\n");
if(pixels_9_7!==16'h083d) $display("ERROR! at (9,7)\n");
if(pixels_10_7!==16'h0285) $display("ERROR! at (10,7)\n");
if(pixels_11_7!==16'h004a) $display("ERROR! at (11,7)\n");
if(pixels_12_7!==16'hfc6a) $display("ERROR! at (12,7)\n");
if(pixels_13_7!==16'hfd5d) $display("ERROR! at (13,7)\n");
if(pixels_14_7!==16'h010e) $display("ERROR! at (14,7)\n");
if(pixels_15_7!==16'h0626) $display("ERROR! at (15,7)\n");
if(pixels_16_7!==16'hfb1c) $display("ERROR! at (16,7)\n");
if(pixels_17_7!==16'h0549) $display("ERROR! at (17,7)\n");
if(pixels_18_7!==16'h00dd) $display("ERROR! at (18,7)\n");
if(pixels_19_7!==16'hf5bc) $display("ERROR! at (19,7)\n");
if(pixels_20_7!==16'h0288) $display("ERROR! at (20,7)\n");
if(pixels_21_7!==16'hf9cc) $display("ERROR! at (21,7)\n");
if(pixels_22_7!==16'hfd19) $display("ERROR! at (22,7)\n");
if(pixels_23_7!==16'hfa2e) $display("ERROR! at (23,7)\n");
if(pixels_24_7!==16'hff93) $display("ERROR! at (24,7)\n");
if(pixels_25_7!==16'hfd8b) $display("ERROR! at (25,7)\n");
if(pixels_26_7!==16'h0032) $display("ERROR! at (26,7)\n");
if(pixels_27_7!==16'hf9f8) $display("ERROR! at (27,7)\n");
if(pixels_28_7!==16'h0026) $display("ERROR! at (28,7)\n");
if(pixels_29_7!==16'h00e9) $display("ERROR! at (29,7)\n");
if(pixels_30_7!==16'hfc3b) $display("ERROR! at (30,7)\n");
if(pixels_31_7!==16'hfcf1) $display("ERROR! at (31,7)\n");
if(pixels_0_8!==16'hff9a) $display("ERROR! at (0,8)\n");
if(pixels_1_8!==16'hfc6f) $display("ERROR! at (1,8)\n");
if(pixels_2_8!==16'hfcf4) $display("ERROR! at (2,8)\n");
if(pixels_3_8!==16'hfc6e) $display("ERROR! at (3,8)\n");
if(pixels_4_8!==16'hfac6) $display("ERROR! at (4,8)\n");
if(pixels_5_8!==16'h068c) $display("ERROR! at (5,8)\n");
if(pixels_6_8!==16'hfc8b) $display("ERROR! at (6,8)\n");
if(pixels_7_8!==16'h0a86) $display("ERROR! at (7,8)\n");
if(pixels_8_8!==16'hf2e8) $display("ERROR! at (8,8)\n");
if(pixels_9_8!==16'h0306) $display("ERROR! at (9,8)\n");
if(pixels_10_8!==16'hf53f) $display("ERROR! at (10,8)\n");
if(pixels_11_8!==16'hfc68) $display("ERROR! at (11,8)\n");
if(pixels_12_8!==16'h0338) $display("ERROR! at (12,8)\n");
if(pixels_13_8!==16'hfb3d) $display("ERROR! at (13,8)\n");
if(pixels_14_8!==16'hfaea) $display("ERROR! at (14,8)\n");
if(pixels_15_8!==16'hfd48) $display("ERROR! at (15,8)\n");
if(pixels_16_8!==16'h00ee) $display("ERROR! at (16,8)\n");
if(pixels_17_8!==16'hfa85) $display("ERROR! at (17,8)\n");
if(pixels_18_8!==16'h022c) $display("ERROR! at (18,8)\n");
if(pixels_19_8!==16'hff3e) $display("ERROR! at (19,8)\n");
if(pixels_20_8!==16'hff83) $display("ERROR! at (20,8)\n");
if(pixels_21_8!==16'h002c) $display("ERROR! at (21,8)\n");
if(pixels_22_8!==16'hfc27) $display("ERROR! at (22,8)\n");
if(pixels_23_8!==16'hfc61) $display("ERROR! at (23,8)\n");
if(pixels_24_8!==16'hf563) $display("ERROR! at (24,8)\n");
if(pixels_25_8!==16'hfc5a) $display("ERROR! at (25,8)\n");
if(pixels_26_8!==16'hfc7b) $display("ERROR! at (26,8)\n");
if(pixels_27_8!==16'h028e) $display("ERROR! at (27,8)\n");
if(pixels_28_8!==16'hf833) $display("ERROR! at (28,8)\n");
if(pixels_29_8!==16'hff58) $display("ERROR! at (29,8)\n");
if(pixels_30_8!==16'hff7a) $display("ERROR! at (30,8)\n");
if(pixels_31_8!==16'h00bb) $display("ERROR! at (31,8)\n");
if(pixels_0_9!==16'h00c8) $display("ERROR! at (0,9)\n");
if(pixels_1_9!==16'h02c5) $display("ERROR! at (1,9)\n");
if(pixels_2_9!==16'hfe23) $display("ERROR! at (2,9)\n");
if(pixels_3_9!==16'h0611) $display("ERROR! at (3,9)\n");
if(pixels_4_9!==16'h0521) $display("ERROR! at (4,9)\n");
if(pixels_5_9!==16'hfcf2) $display("ERROR! at (5,9)\n");
if(pixels_6_9!==16'hffdb) $display("ERROR! at (6,9)\n");
if(pixels_7_9!==16'hfccb) $display("ERROR! at (7,9)\n");
if(pixels_8_9!==16'h009c) $display("ERROR! at (8,9)\n");
if(pixels_9_9!==16'hf28e) $display("ERROR! at (9,9)\n");
if(pixels_10_9!==16'h04c9) $display("ERROR! at (10,9)\n");
if(pixels_11_9!==16'hfaed) $display("ERROR! at (11,9)\n");
if(pixels_12_9!==16'h001c) $display("ERROR! at (12,9)\n");
if(pixels_13_9!==16'hfd3e) $display("ERROR! at (13,9)\n");
if(pixels_14_9!==16'h012d) $display("ERROR! at (14,9)\n");
if(pixels_15_9!==16'h01ad) $display("ERROR! at (15,9)\n");
if(pixels_16_9!==16'h0263) $display("ERROR! at (16,9)\n");
if(pixels_17_9!==16'h035e) $display("ERROR! at (17,9)\n");
if(pixels_18_9!==16'hfff3) $display("ERROR! at (18,9)\n");
if(pixels_19_9!==16'hfab4) $display("ERROR! at (19,9)\n");
if(pixels_20_9!==16'hf455) $display("ERROR! at (20,9)\n");
if(pixels_21_9!==16'hfa51) $display("ERROR! at (21,9)\n");
if(pixels_22_9!==16'hfc98) $display("ERROR! at (22,9)\n");
if(pixels_23_9!==16'hfcba) $display("ERROR! at (23,9)\n");
if(pixels_24_9!==16'h0536) $display("ERROR! at (24,9)\n");
if(pixels_25_9!==16'h0671) $display("ERROR! at (25,9)\n");
if(pixels_26_9!==16'hfdcc) $display("ERROR! at (26,9)\n");
if(pixels_27_9!==16'hfbde) $display("ERROR! at (27,9)\n");
if(pixels_28_9!==16'hfb20) $display("ERROR! at (28,9)\n");
if(pixels_29_9!==16'hfc57) $display("ERROR! at (29,9)\n");
if(pixels_30_9!==16'h0326) $display("ERROR! at (30,9)\n");
if(pixels_31_9!==16'hfe20) $display("ERROR! at (31,9)\n");
if(pixels_0_10!==16'hfefe) $display("ERROR! at (0,10)\n");
if(pixels_1_10!==16'hfe13) $display("ERROR! at (1,10)\n");
if(pixels_2_10!==16'hfa8e) $display("ERROR! at (2,10)\n");
if(pixels_3_10!==16'h0006) $display("ERROR! at (3,10)\n");
if(pixels_4_10!==16'h04f0) $display("ERROR! at (4,10)\n");
if(pixels_5_10!==16'hff6b) $display("ERROR! at (5,10)\n");
if(pixels_6_10!==16'h0630) $display("ERROR! at (6,10)\n");
if(pixels_7_10!==16'h00ee) $display("ERROR! at (7,10)\n");
if(pixels_8_10!==16'hfedc) $display("ERROR! at (8,10)\n");
if(pixels_9_10!==16'hf922) $display("ERROR! at (9,10)\n");
if(pixels_10_10!==16'hfab3) $display("ERROR! at (10,10)\n");
if(pixels_11_10!==16'hf7f5) $display("ERROR! at (11,10)\n");
if(pixels_12_10!==16'hfb43) $display("ERROR! at (12,10)\n");
if(pixels_13_10!==16'hfb7d) $display("ERROR! at (13,10)\n");
if(pixels_14_10!==16'hf97b) $display("ERROR! at (14,10)\n");
if(pixels_15_10!==16'hffda) $display("ERROR! at (15,10)\n");
if(pixels_16_10!==16'h029c) $display("ERROR! at (16,10)\n");
if(pixels_17_10!==16'hfdd4) $display("ERROR! at (17,10)\n");
if(pixels_18_10!==16'hfd4e) $display("ERROR! at (18,10)\n");
if(pixels_19_10!==16'hfdb3) $display("ERROR! at (19,10)\n");
if(pixels_20_10!==16'hfc12) $display("ERROR! at (20,10)\n");
if(pixels_21_10!==16'h0141) $display("ERROR! at (21,10)\n");
if(pixels_22_10!==16'h0492) $display("ERROR! at (22,10)\n");
if(pixels_23_10!==16'hf9a2) $display("ERROR! at (23,10)\n");
if(pixels_24_10!==16'hf920) $display("ERROR! at (24,10)\n");
if(pixels_25_10!==16'hfbfe) $display("ERROR! at (25,10)\n");
if(pixels_26_10!==16'h007c) $display("ERROR! at (26,10)\n");
if(pixels_27_10!==16'h00d1) $display("ERROR! at (27,10)\n");
if(pixels_28_10!==16'h0375) $display("ERROR! at (28,10)\n");
if(pixels_29_10!==16'hfc0c) $display("ERROR! at (29,10)\n");
if(pixels_30_10!==16'hfdf6) $display("ERROR! at (30,10)\n");
if(pixels_31_10!==16'hfed3) $display("ERROR! at (31,10)\n");
if(pixels_0_11!==16'h00d2) $display("ERROR! at (0,11)\n");
if(pixels_1_11!==16'h049d) $display("ERROR! at (1,11)\n");
if(pixels_2_11!==16'h0151) $display("ERROR! at (2,11)\n");
if(pixels_3_11!==16'hfd96) $display("ERROR! at (3,11)\n");
if(pixels_4_11!==16'h0302) $display("ERROR! at (4,11)\n");
if(pixels_5_11!==16'hfbc9) $display("ERROR! at (5,11)\n");
if(pixels_6_11!==16'hfb36) $display("ERROR! at (6,11)\n");
if(pixels_7_11!==16'h0220) $display("ERROR! at (7,11)\n");
if(pixels_8_11!==16'h0049) $display("ERROR! at (8,11)\n");
if(pixels_9_11!==16'h025a) $display("ERROR! at (9,11)\n");
if(pixels_10_11!==16'hff7a) $display("ERROR! at (10,11)\n");
if(pixels_11_11!==16'h0383) $display("ERROR! at (11,11)\n");
if(pixels_12_11!==16'h0076) $display("ERROR! at (12,11)\n");
if(pixels_13_11!==16'h028b) $display("ERROR! at (13,11)\n");
if(pixels_14_11!==16'hffbe) $display("ERROR! at (14,11)\n");
if(pixels_15_11!==16'hff1b) $display("ERROR! at (15,11)\n");
if(pixels_16_11!==16'hfd9c) $display("ERROR! at (16,11)\n");
if(pixels_17_11!==16'hff62) $display("ERROR! at (17,11)\n");
if(pixels_18_11!==16'hff48) $display("ERROR! at (18,11)\n");
if(pixels_19_11!==16'hf72f) $display("ERROR! at (19,11)\n");
if(pixels_20_11!==16'hfc90) $display("ERROR! at (20,11)\n");
if(pixels_21_11!==16'hfbbc) $display("ERROR! at (21,11)\n");
if(pixels_22_11!==16'hfeb7) $display("ERROR! at (22,11)\n");
if(pixels_23_11!==16'h0338) $display("ERROR! at (23,11)\n");
if(pixels_24_11!==16'h0231) $display("ERROR! at (24,11)\n");
if(pixels_25_11!==16'h0779) $display("ERROR! at (25,11)\n");
if(pixels_26_11!==16'h0559) $display("ERROR! at (26,11)\n");
if(pixels_27_11!==16'hff43) $display("ERROR! at (27,11)\n");
if(pixels_28_11!==16'h00a6) $display("ERROR! at (28,11)\n");
if(pixels_29_11!==16'h007b) $display("ERROR! at (29,11)\n");
if(pixels_30_11!==16'h0159) $display("ERROR! at (30,11)\n");
if(pixels_31_11!==16'h01c1) $display("ERROR! at (31,11)\n");
if(pixels_0_12!==16'hff19) $display("ERROR! at (0,12)\n");
if(pixels_1_12!==16'hfe6a) $display("ERROR! at (1,12)\n");
if(pixels_2_12!==16'hfcd7) $display("ERROR! at (2,12)\n");
if(pixels_3_12!==16'hff17) $display("ERROR! at (3,12)\n");
if(pixels_4_12!==16'h04c3) $display("ERROR! at (4,12)\n");
if(pixels_5_12!==16'h0541) $display("ERROR! at (5,12)\n");
if(pixels_6_12!==16'hfa25) $display("ERROR! at (6,12)\n");
if(pixels_7_12!==16'hf9e0) $display("ERROR! at (7,12)\n");
if(pixels_8_12!==16'hfc99) $display("ERROR! at (8,12)\n");
if(pixels_9_12!==16'hf423) $display("ERROR! at (9,12)\n");
if(pixels_10_12!==16'h00e7) $display("ERROR! at (10,12)\n");
if(pixels_11_12!==16'hfabd) $display("ERROR! at (11,12)\n");
if(pixels_12_12!==16'h07e2) $display("ERROR! at (12,12)\n");
if(pixels_13_12!==16'hffc8) $display("ERROR! at (13,12)\n");
if(pixels_14_12!==16'h0026) $display("ERROR! at (14,12)\n");
if(pixels_15_12!==16'hf772) $display("ERROR! at (15,12)\n");
if(pixels_16_12!==16'h0051) $display("ERROR! at (16,12)\n");
if(pixels_17_12!==16'hff61) $display("ERROR! at (17,12)\n");
if(pixels_18_12!==16'hfe4a) $display("ERROR! at (18,12)\n");
if(pixels_19_12!==16'hfad6) $display("ERROR! at (19,12)\n");
if(pixels_20_12!==16'hffa5) $display("ERROR! at (20,12)\n");
if(pixels_21_12!==16'hfe16) $display("ERROR! at (21,12)\n");
if(pixels_22_12!==16'h026f) $display("ERROR! at (22,12)\n");
if(pixels_23_12!==16'h01fa) $display("ERROR! at (23,12)\n");
if(pixels_24_12!==16'h00ac) $display("ERROR! at (24,12)\n");
if(pixels_25_12!==16'hf69a) $display("ERROR! at (25,12)\n");
if(pixels_26_12!==16'h0557) $display("ERROR! at (26,12)\n");
if(pixels_27_12!==16'h0464) $display("ERROR! at (27,12)\n");
if(pixels_28_12!==16'h0320) $display("ERROR! at (28,12)\n");
if(pixels_29_12!==16'h029e) $display("ERROR! at (29,12)\n");
if(pixels_30_12!==16'hff8d) $display("ERROR! at (30,12)\n");
if(pixels_31_12!==16'hff52) $display("ERROR! at (31,12)\n");
if(pixels_0_13!==16'h00fe) $display("ERROR! at (0,13)\n");
if(pixels_1_13!==16'hfccb) $display("ERROR! at (1,13)\n");
if(pixels_2_13!==16'h07d4) $display("ERROR! at (2,13)\n");
if(pixels_3_13!==16'hfcfc) $display("ERROR! at (3,13)\n");
if(pixels_4_13!==16'hfdab) $display("ERROR! at (4,13)\n");
if(pixels_5_13!==16'h05e1) $display("ERROR! at (5,13)\n");
if(pixels_6_13!==16'h03e1) $display("ERROR! at (6,13)\n");
if(pixels_7_13!==16'hf972) $display("ERROR! at (7,13)\n");
if(pixels_8_13!==16'h0471) $display("ERROR! at (8,13)\n");
if(pixels_9_13!==16'hfde4) $display("ERROR! at (9,13)\n");
if(pixels_10_13!==16'h0586) $display("ERROR! at (10,13)\n");
if(pixels_11_13!==16'h00e1) $display("ERROR! at (11,13)\n");
if(pixels_12_13!==16'hfd5e) $display("ERROR! at (12,13)\n");
if(pixels_13_13!==16'h000e) $display("ERROR! at (13,13)\n");
if(pixels_14_13!==16'h04d1) $display("ERROR! at (14,13)\n");
if(pixels_15_13!==16'hfe79) $display("ERROR! at (15,13)\n");
if(pixels_16_13!==16'hfa4e) $display("ERROR! at (16,13)\n");
if(pixels_17_13!==16'hfd56) $display("ERROR! at (17,13)\n");
if(pixels_18_13!==16'hfd5a) $display("ERROR! at (18,13)\n");
if(pixels_19_13!==16'hfe8e) $display("ERROR! at (19,13)\n");
if(pixels_20_13!==16'hf714) $display("ERROR! at (20,13)\n");
if(pixels_21_13!==16'h0790) $display("ERROR! at (21,13)\n");
if(pixels_22_13!==16'hfe35) $display("ERROR! at (22,13)\n");
if(pixels_23_13!==16'h02a7) $display("ERROR! at (23,13)\n");
if(pixels_24_13!==16'hfaac) $display("ERROR! at (24,13)\n");
if(pixels_25_13!==16'h0590) $display("ERROR! at (25,13)\n");
if(pixels_26_13!==16'hffe3) $display("ERROR! at (26,13)\n");
if(pixels_27_13!==16'h080a) $display("ERROR! at (27,13)\n");
if(pixels_28_13!==16'hfe10) $display("ERROR! at (28,13)\n");
if(pixels_29_13!==16'hff48) $display("ERROR! at (29,13)\n");
if(pixels_30_13!==16'hff27) $display("ERROR! at (30,13)\n");
if(pixels_31_13!==16'hfeb1) $display("ERROR! at (31,13)\n");
if(pixels_0_14!==16'hfd2c) $display("ERROR! at (0,14)\n");
if(pixels_1_14!==16'h002c) $display("ERROR! at (1,14)\n");
if(pixels_2_14!==16'hfde4) $display("ERROR! at (2,14)\n");
if(pixels_3_14!==16'h0436) $display("ERROR! at (3,14)\n");
if(pixels_4_14!==16'hfd50) $display("ERROR! at (4,14)\n");
if(pixels_5_14!==16'h0109) $display("ERROR! at (5,14)\n");
if(pixels_6_14!==16'h033e) $display("ERROR! at (6,14)\n");
if(pixels_7_14!==16'hfea6) $display("ERROR! at (7,14)\n");
if(pixels_8_14!==16'h05e2) $display("ERROR! at (8,14)\n");
if(pixels_9_14!==16'hfe7e) $display("ERROR! at (9,14)\n");
if(pixels_10_14!==16'hfc34) $display("ERROR! at (10,14)\n");
if(pixels_11_14!==16'h014a) $display("ERROR! at (11,14)\n");
if(pixels_12_14!==16'hffe3) $display("ERROR! at (12,14)\n");
if(pixels_13_14!==16'h03dd) $display("ERROR! at (13,14)\n");
if(pixels_14_14!==16'h0662) $display("ERROR! at (14,14)\n");
if(pixels_15_14!==16'hfc84) $display("ERROR! at (15,14)\n");
if(pixels_16_14!==16'h0173) $display("ERROR! at (16,14)\n");
if(pixels_17_14!==16'h04d7) $display("ERROR! at (17,14)\n");
if(pixels_18_14!==16'h04d2) $display("ERROR! at (18,14)\n");
if(pixels_19_14!==16'hff51) $display("ERROR! at (19,14)\n");
if(pixels_20_14!==16'h0263) $display("ERROR! at (20,14)\n");
if(pixels_21_14!==16'h0093) $display("ERROR! at (21,14)\n");
if(pixels_22_14!==16'h074f) $display("ERROR! at (22,14)\n");
if(pixels_23_14!==16'h024b) $display("ERROR! at (23,14)\n");
if(pixels_24_14!==16'h02dc) $display("ERROR! at (24,14)\n");
if(pixels_25_14!==16'hfcb3) $display("ERROR! at (25,14)\n");
if(pixels_26_14!==16'h0215) $display("ERROR! at (26,14)\n");
if(pixels_27_14!==16'h00a9) $display("ERROR! at (27,14)\n");
if(pixels_28_14!==16'h09fe) $display("ERROR! at (28,14)\n");
if(pixels_29_14!==16'hfda0) $display("ERROR! at (29,14)\n");
if(pixels_30_14!==16'hff15) $display("ERROR! at (30,14)\n");
if(pixels_31_14!==16'hfe7b) $display("ERROR! at (31,14)\n");
if(pixels_0_15!==16'h027d) $display("ERROR! at (0,15)\n");
if(pixels_1_15!==16'hffc3) $display("ERROR! at (1,15)\n");
if(pixels_2_15!==16'h0257) $display("ERROR! at (2,15)\n");
if(pixels_3_15!==16'h04d5) $display("ERROR! at (3,15)\n");
if(pixels_4_15!==16'h0b5f) $display("ERROR! at (4,15)\n");
if(pixels_5_15!==16'hfe42) $display("ERROR! at (5,15)\n");
if(pixels_6_15!==16'h05c2) $display("ERROR! at (6,15)\n");
if(pixels_7_15!==16'h03e2) $display("ERROR! at (7,15)\n");
if(pixels_8_15!==16'hfc37) $display("ERROR! at (8,15)\n");
if(pixels_9_15!==16'h046c) $display("ERROR! at (9,15)\n");
if(pixels_10_15!==16'h00c0) $display("ERROR! at (10,15)\n");
if(pixels_11_15!==16'hff28) $display("ERROR! at (11,15)\n");
if(pixels_12_15!==16'h01e0) $display("ERROR! at (12,15)\n");
if(pixels_13_15!==16'hf2e9) $display("ERROR! at (13,15)\n");
if(pixels_14_15!==16'h0338) $display("ERROR! at (14,15)\n");
if(pixels_15_15!==16'hfe24) $display("ERROR! at (15,15)\n");
if(pixels_16_15!==16'hfc8e) $display("ERROR! at (16,15)\n");
if(pixels_17_15!==16'hfb52) $display("ERROR! at (17,15)\n");
if(pixels_18_15!==16'h002f) $display("ERROR! at (18,15)\n");
if(pixels_19_15!==16'h037b) $display("ERROR! at (19,15)\n");
if(pixels_20_15!==16'h039e) $display("ERROR! at (20,15)\n");
if(pixels_21_15!==16'hff0b) $display("ERROR! at (21,15)\n");
if(pixels_22_15!==16'h010f) $display("ERROR! at (22,15)\n");
if(pixels_23_15!==16'h0194) $display("ERROR! at (23,15)\n");
if(pixels_24_15!==16'h0042) $display("ERROR! at (24,15)\n");
if(pixels_25_15!==16'hff4a) $display("ERROR! at (25,15)\n");
if(pixels_26_15!==16'h07a1) $display("ERROR! at (26,15)\n");
if(pixels_27_15!==16'h0765) $display("ERROR! at (27,15)\n");
if(pixels_28_15!==16'h00f2) $display("ERROR! at (28,15)\n");
if(pixels_29_15!==16'hfdaf) $display("ERROR! at (29,15)\n");
if(pixels_30_15!==16'hfd85) $display("ERROR! at (30,15)\n");
if(pixels_31_15!==16'hfe94) $display("ERROR! at (31,15)\n");
if(pixels_0_16!==16'hfe8e) $display("ERROR! at (0,16)\n");
if(pixels_1_16!==16'hfe7e) $display("ERROR! at (1,16)\n");
if(pixels_2_16!==16'hfe22) $display("ERROR! at (2,16)\n");
if(pixels_3_16!==16'h0093) $display("ERROR! at (3,16)\n");
if(pixels_4_16!==16'h0376) $display("ERROR! at (4,16)\n");
if(pixels_5_16!==16'h0501) $display("ERROR! at (5,16)\n");
if(pixels_6_16!==16'hfee8) $display("ERROR! at (6,16)\n");
if(pixels_7_16!==16'h00e4) $display("ERROR! at (7,16)\n");
if(pixels_8_16!==16'h05e7) $display("ERROR! at (8,16)\n");
if(pixels_9_16!==16'h04c5) $display("ERROR! at (9,16)\n");
if(pixels_10_16!==16'h0297) $display("ERROR! at (10,16)\n");
if(pixels_11_16!==16'hf616) $display("ERROR! at (11,16)\n");
if(pixels_12_16!==16'h0404) $display("ERROR! at (12,16)\n");
if(pixels_13_16!==16'h04ec) $display("ERROR! at (13,16)\n");
if(pixels_14_16!==16'h0388) $display("ERROR! at (14,16)\n");
if(pixels_15_16!==16'h09bd) $display("ERROR! at (15,16)\n");
if(pixels_16_16!==16'h00fe) $display("ERROR! at (16,16)\n");
if(pixels_17_16!==16'h091e) $display("ERROR! at (17,16)\n");
if(pixels_18_16!==16'h0325) $display("ERROR! at (18,16)\n");
if(pixels_19_16!==16'h03e7) $display("ERROR! at (19,16)\n");
if(pixels_20_16!==16'hfd88) $display("ERROR! at (20,16)\n");
if(pixels_21_16!==16'h01b5) $display("ERROR! at (21,16)\n");
if(pixels_22_16!==16'hfaf5) $display("ERROR! at (22,16)\n");
if(pixels_23_16!==16'h00c0) $display("ERROR! at (23,16)\n");
if(pixels_24_16!==16'hf766) $display("ERROR! at (24,16)\n");
if(pixels_25_16!==16'h0734) $display("ERROR! at (25,16)\n");
if(pixels_26_16!==16'hff08) $display("ERROR! at (26,16)\n");
if(pixels_27_16!==16'h04fb) $display("ERROR! at (27,16)\n");
if(pixels_28_16!==16'hfbd3) $display("ERROR! at (28,16)\n");
if(pixels_29_16!==16'h0060) $display("ERROR! at (29,16)\n");
if(pixels_30_16!==16'hfc4d) $display("ERROR! at (30,16)\n");
if(pixels_31_16!==16'hff19) $display("ERROR! at (31,16)\n");
if(pixels_0_17!==16'h013e) $display("ERROR! at (0,17)\n");
if(pixels_1_17!==16'hff37) $display("ERROR! at (1,17)\n");
if(pixels_2_17!==16'hfff2) $display("ERROR! at (2,17)\n");
if(pixels_3_17!==16'h00a5) $display("ERROR! at (3,17)\n");
if(pixels_4_17!==16'hfd7c) $display("ERROR! at (4,17)\n");
if(pixels_5_17!==16'h00e5) $display("ERROR! at (5,17)\n");
if(pixels_6_17!==16'h05c4) $display("ERROR! at (6,17)\n");
if(pixels_7_17!==16'hff95) $display("ERROR! at (7,17)\n");
if(pixels_8_17!==16'h006a) $display("ERROR! at (8,17)\n");
if(pixels_9_17!==16'hfe74) $display("ERROR! at (9,17)\n");
if(pixels_10_17!==16'h014b) $display("ERROR! at (10,17)\n");
if(pixels_11_17!==16'h06ec) $display("ERROR! at (11,17)\n");
if(pixels_12_17!==16'hff8a) $display("ERROR! at (12,17)\n");
if(pixels_13_17!==16'h03c8) $display("ERROR! at (13,17)\n");
if(pixels_14_17!==16'hf397) $display("ERROR! at (14,17)\n");
if(pixels_15_17!==16'h00bc) $display("ERROR! at (15,17)\n");
if(pixels_16_17!==16'h06ab) $display("ERROR! at (16,17)\n");
if(pixels_17_17!==16'h002c) $display("ERROR! at (17,17)\n");
if(pixels_18_17!==16'h02a6) $display("ERROR! at (18,17)\n");
if(pixels_19_17!==16'h0310) $display("ERROR! at (19,17)\n");
if(pixels_20_17!==16'h0041) $display("ERROR! at (20,17)\n");
if(pixels_21_17!==16'h01b1) $display("ERROR! at (21,17)\n");
if(pixels_22_17!==16'hff8d) $display("ERROR! at (22,17)\n");
if(pixels_23_17!==16'h0097) $display("ERROR! at (23,17)\n");
if(pixels_24_17!==16'h05b2) $display("ERROR! at (24,17)\n");
if(pixels_25_17!==16'hff1f) $display("ERROR! at (25,17)\n");
if(pixels_26_17!==16'hfcfa) $display("ERROR! at (26,17)\n");
if(pixels_27_17!==16'hff53) $display("ERROR! at (27,17)\n");
if(pixels_28_17!==16'h008b) $display("ERROR! at (28,17)\n");
if(pixels_29_17!==16'hfe07) $display("ERROR! at (29,17)\n");
if(pixels_30_17!==16'hfc4c) $display("ERROR! at (30,17)\n");
if(pixels_31_17!==16'h0083) $display("ERROR! at (31,17)\n");
if(pixels_0_18!==16'h0241) $display("ERROR! at (0,18)\n");
if(pixels_1_18!==16'hfb55) $display("ERROR! at (1,18)\n");
if(pixels_2_18!==16'h0075) $display("ERROR! at (2,18)\n");
if(pixels_3_18!==16'h04dc) $display("ERROR! at (3,18)\n");
if(pixels_4_18!==16'hfd4c) $display("ERROR! at (4,18)\n");
if(pixels_5_18!==16'h032f) $display("ERROR! at (5,18)\n");
if(pixels_6_18!==16'h0275) $display("ERROR! at (6,18)\n");
if(pixels_7_18!==16'h01d5) $display("ERROR! at (7,18)\n");
if(pixels_8_18!==16'hfdf9) $display("ERROR! at (8,18)\n");
if(pixels_9_18!==16'h0975) $display("ERROR! at (9,18)\n");
if(pixels_10_18!==16'hfef0) $display("ERROR! at (10,18)\n");
if(pixels_11_18!==16'h0044) $display("ERROR! at (11,18)\n");
if(pixels_12_18!==16'h01fb) $display("ERROR! at (12,18)\n");
if(pixels_13_18!==16'hffe7) $display("ERROR! at (13,18)\n");
if(pixels_14_18!==16'h03e5) $display("ERROR! at (14,18)\n");
if(pixels_15_18!==16'hfda2) $display("ERROR! at (15,18)\n");
if(pixels_16_18!==16'h0369) $display("ERROR! at (16,18)\n");
if(pixels_17_18!==16'hfd18) $display("ERROR! at (17,18)\n");
if(pixels_18_18!==16'hfbf7) $display("ERROR! at (18,18)\n");
if(pixels_19_18!==16'hffa5) $display("ERROR! at (19,18)\n");
if(pixels_20_18!==16'h0034) $display("ERROR! at (20,18)\n");
if(pixels_21_18!==16'h02ff) $display("ERROR! at (21,18)\n");
if(pixels_22_18!==16'hfeec) $display("ERROR! at (22,18)\n");
if(pixels_23_18!==16'hfe71) $display("ERROR! at (23,18)\n");
if(pixels_24_18!==16'h0092) $display("ERROR! at (24,18)\n");
if(pixels_25_18!==16'h0328) $display("ERROR! at (25,18)\n");
if(pixels_26_18!==16'h03d2) $display("ERROR! at (26,18)\n");
if(pixels_27_18!==16'h068e) $display("ERROR! at (27,18)\n");
if(pixels_28_18!==16'hfe9e) $display("ERROR! at (28,18)\n");
if(pixels_29_18!==16'hfdea) $display("ERROR! at (29,18)\n");
if(pixels_30_18!==16'h0660) $display("ERROR! at (30,18)\n");
if(pixels_31_18!==16'h0148) $display("ERROR! at (31,18)\n");
if(pixels_0_19!==16'hfe49) $display("ERROR! at (0,19)\n");
if(pixels_1_19!==16'h0064) $display("ERROR! at (1,19)\n");
if(pixels_2_19!==16'hfe48) $display("ERROR! at (2,19)\n");
if(pixels_3_19!==16'h022a) $display("ERROR! at (3,19)\n");
if(pixels_4_19!==16'h076e) $display("ERROR! at (4,19)\n");
if(pixels_5_19!==16'h017d) $display("ERROR! at (5,19)\n");
if(pixels_6_19!==16'hfe07) $display("ERROR! at (6,19)\n");
if(pixels_7_19!==16'h01ea) $display("ERROR! at (7,19)\n");
if(pixels_8_19!==16'hfcdf) $display("ERROR! at (8,19)\n");
if(pixels_9_19!==16'hfdb9) $display("ERROR! at (9,19)\n");
if(pixels_10_19!==16'h001c) $display("ERROR! at (10,19)\n");
if(pixels_11_19!==16'hfc0d) $display("ERROR! at (11,19)\n");
if(pixels_12_19!==16'h07c9) $display("ERROR! at (12,19)\n");
if(pixels_13_19!==16'h0092) $display("ERROR! at (13,19)\n");
if(pixels_14_19!==16'h0278) $display("ERROR! at (14,19)\n");
if(pixels_15_19!==16'h01c3) $display("ERROR! at (15,19)\n");
if(pixels_16_19!==16'h00fe) $display("ERROR! at (16,19)\n");
if(pixels_17_19!==16'h0719) $display("ERROR! at (17,19)\n");
if(pixels_18_19!==16'hfda8) $display("ERROR! at (18,19)\n");
if(pixels_19_19!==16'hfefa) $display("ERROR! at (19,19)\n");
if(pixels_20_19!==16'h04d1) $display("ERROR! at (20,19)\n");
if(pixels_21_19!==16'h0191) $display("ERROR! at (21,19)\n");
if(pixels_22_19!==16'hff2b) $display("ERROR! at (22,19)\n");
if(pixels_23_19!==16'h026d) $display("ERROR! at (23,19)\n");
if(pixels_24_19!==16'hfa72) $display("ERROR! at (24,19)\n");
if(pixels_25_19!==16'h0646) $display("ERROR! at (25,19)\n");
if(pixels_26_19!==16'hfb69) $display("ERROR! at (26,19)\n");
if(pixels_27_19!==16'hfb04) $display("ERROR! at (27,19)\n");
if(pixels_28_19!==16'hff6e) $display("ERROR! at (28,19)\n");
if(pixels_29_19!==16'h02ef) $display("ERROR! at (29,19)\n");
if(pixels_30_19!==16'hffd1) $display("ERROR! at (30,19)\n");
if(pixels_31_19!==16'h000f) $display("ERROR! at (31,19)\n");
if(pixels_0_20!==16'h0332) $display("ERROR! at (0,20)\n");
if(pixels_1_20!==16'h01e6) $display("ERROR! at (1,20)\n");
if(pixels_2_20!==16'hfd7e) $display("ERROR! at (2,20)\n");
if(pixels_3_20!==16'h00f2) $display("ERROR! at (3,20)\n");
if(pixels_4_20!==16'h025f) $display("ERROR! at (4,20)\n");
if(pixels_5_20!==16'hff8d) $display("ERROR! at (5,20)\n");
if(pixels_6_20!==16'hfd4e) $display("ERROR! at (6,20)\n");
if(pixels_7_20!==16'h04a2) $display("ERROR! at (7,20)\n");
if(pixels_8_20!==16'hfc7e) $display("ERROR! at (8,20)\n");
if(pixels_9_20!==16'hfeac) $display("ERROR! at (9,20)\n");
if(pixels_10_20!==16'h021c) $display("ERROR! at (10,20)\n");
if(pixels_11_20!==16'hff64) $display("ERROR! at (11,20)\n");
if(pixels_12_20!==16'hfa17) $display("ERROR! at (12,20)\n");
if(pixels_13_20!==16'h041c) $display("ERROR! at (13,20)\n");
if(pixels_14_20!==16'hfa4a) $display("ERROR! at (14,20)\n");
if(pixels_15_20!==16'h01c3) $display("ERROR! at (15,20)\n");
if(pixels_16_20!==16'hfac1) $display("ERROR! at (16,20)\n");
if(pixels_17_20!==16'h03e0) $display("ERROR! at (17,20)\n");
if(pixels_18_20!==16'hfe03) $display("ERROR! at (18,20)\n");
if(pixels_19_20!==16'hf6d6) $display("ERROR! at (19,20)\n");
if(pixels_20_20!==16'hfa5a) $display("ERROR! at (20,20)\n");
if(pixels_21_20!==16'hfbf7) $display("ERROR! at (21,20)\n");
if(pixels_22_20!==16'hfc2f) $display("ERROR! at (22,20)\n");
if(pixels_23_20!==16'h04ba) $display("ERROR! at (23,20)\n");
if(pixels_24_20!==16'h0480) $display("ERROR! at (24,20)\n");
if(pixels_25_20!==16'hff4b) $display("ERROR! at (25,20)\n");
if(pixels_26_20!==16'hff12) $display("ERROR! at (26,20)\n");
if(pixels_27_20!==16'h0390) $display("ERROR! at (27,20)\n");
if(pixels_28_20!==16'h01e1) $display("ERROR! at (28,20)\n");
if(pixels_29_20!==16'h014a) $display("ERROR! at (29,20)\n");
if(pixels_30_20!==16'hffe3) $display("ERROR! at (30,20)\n");
if(pixels_31_20!==16'h03f9) $display("ERROR! at (31,20)\n");
if(pixels_0_21!==16'hffc7) $display("ERROR! at (0,21)\n");
if(pixels_1_21!==16'h02e6) $display("ERROR! at (1,21)\n");
if(pixels_2_21!==16'h0327) $display("ERROR! at (2,21)\n");
if(pixels_3_21!==16'hfe35) $display("ERROR! at (3,21)\n");
if(pixels_4_21!==16'h05e4) $display("ERROR! at (4,21)\n");
if(pixels_5_21!==16'h01ae) $display("ERROR! at (5,21)\n");
if(pixels_6_21!==16'h019a) $display("ERROR! at (6,21)\n");
if(pixels_7_21!==16'hfe38) $display("ERROR! at (7,21)\n");
if(pixels_8_21!==16'hfcbb) $display("ERROR! at (8,21)\n");
if(pixels_9_21!==16'hfe9e) $display("ERROR! at (9,21)\n");
if(pixels_10_21!==16'hfca2) $display("ERROR! at (10,21)\n");
if(pixels_11_21!==16'hfe6f) $display("ERROR! at (11,21)\n");
if(pixels_12_21!==16'hfdbd) $display("ERROR! at (12,21)\n");
if(pixels_13_21!==16'hfeb0) $display("ERROR! at (13,21)\n");
if(pixels_14_21!==16'h033e) $display("ERROR! at (14,21)\n");
if(pixels_15_21!==16'hffd8) $display("ERROR! at (15,21)\n");
if(pixels_16_21!==16'h0497) $display("ERROR! at (16,21)\n");
if(pixels_17_21!==16'hfae8) $display("ERROR! at (17,21)\n");
if(pixels_18_21!==16'hfb35) $display("ERROR! at (18,21)\n");
if(pixels_19_21!==16'hfba5) $display("ERROR! at (19,21)\n");
if(pixels_20_21!==16'hf78e) $display("ERROR! at (20,21)\n");
if(pixels_21_21!==16'h01be) $display("ERROR! at (21,21)\n");
if(pixels_22_21!==16'hf975) $display("ERROR! at (22,21)\n");
if(pixels_23_21!==16'h006b) $display("ERROR! at (23,21)\n");
if(pixels_24_21!==16'hfe5a) $display("ERROR! at (24,21)\n");
if(pixels_25_21!==16'hfead) $display("ERROR! at (25,21)\n");
if(pixels_26_21!==16'hff5d) $display("ERROR! at (26,21)\n");
if(pixels_27_21!==16'h037b) $display("ERROR! at (27,21)\n");
if(pixels_28_21!==16'h00f6) $display("ERROR! at (28,21)\n");
if(pixels_29_21!==16'h03ef) $display("ERROR! at (29,21)\n");
if(pixels_30_21!==16'h08b7) $display("ERROR! at (30,21)\n");
if(pixels_31_21!==16'h0108) $display("ERROR! at (31,21)\n");
if(pixels_0_22!==16'hffb1) $display("ERROR! at (0,22)\n");
if(pixels_1_22!==16'h023f) $display("ERROR! at (1,22)\n");
if(pixels_2_22!==16'hfd92) $display("ERROR! at (2,22)\n");
if(pixels_3_22!==16'hfd97) $display("ERROR! at (3,22)\n");
if(pixels_4_22!==16'hf9a2) $display("ERROR! at (4,22)\n");
if(pixels_5_22!==16'h0692) $display("ERROR! at (5,22)\n");
if(pixels_6_22!==16'hf990) $display("ERROR! at (6,22)\n");
if(pixels_7_22!==16'hfd33) $display("ERROR! at (7,22)\n");
if(pixels_8_22!==16'h010b) $display("ERROR! at (8,22)\n");
if(pixels_9_22!==16'hf80b) $display("ERROR! at (9,22)\n");
if(pixels_10_22!==16'hfe94) $display("ERROR! at (10,22)\n");
if(pixels_11_22!==16'hf807) $display("ERROR! at (11,22)\n");
if(pixels_12_22!==16'hf7bb) $display("ERROR! at (12,22)\n");
if(pixels_13_22!==16'hf98a) $display("ERROR! at (13,22)\n");
if(pixels_14_22!==16'hfdbc) $display("ERROR! at (14,22)\n");
if(pixels_15_22!==16'hfff1) $display("ERROR! at (15,22)\n");
if(pixels_16_22!==16'h0686) $display("ERROR! at (16,22)\n");
if(pixels_17_22!==16'h0216) $display("ERROR! at (17,22)\n");
if(pixels_18_22!==16'hfe09) $display("ERROR! at (18,22)\n");
if(pixels_19_22!==16'h017e) $display("ERROR! at (19,22)\n");
if(pixels_20_22!==16'hfcbd) $display("ERROR! at (20,22)\n");
if(pixels_21_22!==16'hf8a5) $display("ERROR! at (21,22)\n");
if(pixels_22_22!==16'h0286) $display("ERROR! at (22,22)\n");
if(pixels_23_22!==16'hf82c) $display("ERROR! at (23,22)\n");
if(pixels_24_22!==16'hfd98) $display("ERROR! at (24,22)\n");
if(pixels_25_22!==16'h0026) $display("ERROR! at (25,22)\n");
if(pixels_26_22!==16'hfca8) $display("ERROR! at (26,22)\n");
if(pixels_27_22!==16'hf88a) $display("ERROR! at (27,22)\n");
if(pixels_28_22!==16'h013e) $display("ERROR! at (28,22)\n");
if(pixels_29_22!==16'h02f5) $display("ERROR! at (29,22)\n");
if(pixels_30_22!==16'hfead) $display("ERROR! at (30,22)\n");
if(pixels_31_22!==16'hfdb3) $display("ERROR! at (31,22)\n");
if(pixels_0_23!==16'h0072) $display("ERROR! at (0,23)\n");
if(pixels_1_23!==16'hfe3d) $display("ERROR! at (1,23)\n");
if(pixels_2_23!==16'hffd8) $display("ERROR! at (2,23)\n");
if(pixels_3_23!==16'hfef1) $display("ERROR! at (3,23)\n");
if(pixels_4_23!==16'hfcea) $display("ERROR! at (4,23)\n");
if(pixels_5_23!==16'hfc1b) $display("ERROR! at (5,23)\n");
if(pixels_6_23!==16'h0639) $display("ERROR! at (6,23)\n");
if(pixels_7_23!==16'h0091) $display("ERROR! at (7,23)\n");
if(pixels_8_23!==16'hfe67) $display("ERROR! at (8,23)\n");
if(pixels_9_23!==16'h00b1) $display("ERROR! at (9,23)\n");
if(pixels_10_23!==16'hf98c) $display("ERROR! at (10,23)\n");
if(pixels_11_23!==16'hfee5) $display("ERROR! at (11,23)\n");
if(pixels_12_23!==16'h0105) $display("ERROR! at (12,23)\n");
if(pixels_13_23!==16'h0880) $display("ERROR! at (13,23)\n");
if(pixels_14_23!==16'hfd41) $display("ERROR! at (14,23)\n");
if(pixels_15_23!==16'hfb85) $display("ERROR! at (15,23)\n");
if(pixels_16_23!==16'hfbc6) $display("ERROR! at (16,23)\n");
if(pixels_17_23!==16'h05a6) $display("ERROR! at (17,23)\n");
if(pixels_18_23!==16'hfb31) $display("ERROR! at (18,23)\n");
if(pixels_19_23!==16'hfacd) $display("ERROR! at (19,23)\n");
if(pixels_20_23!==16'h0015) $display("ERROR! at (20,23)\n");
if(pixels_21_23!==16'hfc54) $display("ERROR! at (21,23)\n");
if(pixels_22_23!==16'hfe64) $display("ERROR! at (22,23)\n");
if(pixels_23_23!==16'h05e2) $display("ERROR! at (23,23)\n");
if(pixels_24_23!==16'hfd5d) $display("ERROR! at (24,23)\n");
if(pixels_25_23!==16'hfd9b) $display("ERROR! at (25,23)\n");
if(pixels_26_23!==16'hff19) $display("ERROR! at (26,23)\n");
if(pixels_27_23!==16'h021e) $display("ERROR! at (27,23)\n");
if(pixels_28_23!==16'h03af) $display("ERROR! at (28,23)\n");
if(pixels_29_23!==16'h04e8) $display("ERROR! at (29,23)\n");
if(pixels_30_23!==16'hfeac) $display("ERROR! at (30,23)\n");
if(pixels_31_23!==16'h014f) $display("ERROR! at (31,23)\n");
if(pixels_0_24!==16'hff66) $display("ERROR! at (0,24)\n");
if(pixels_1_24!==16'h0060) $display("ERROR! at (1,24)\n");
if(pixels_2_24!==16'h0173) $display("ERROR! at (2,24)\n");
if(pixels_3_24!==16'h0232) $display("ERROR! at (3,24)\n");
if(pixels_4_24!==16'hffaa) $display("ERROR! at (4,24)\n");
if(pixels_5_24!==16'h0684) $display("ERROR! at (5,24)\n");
if(pixels_6_24!==16'hffb9) $display("ERROR! at (6,24)\n");
if(pixels_7_24!==16'hfe21) $display("ERROR! at (7,24)\n");
if(pixels_8_24!==16'hf820) $display("ERROR! at (8,24)\n");
if(pixels_9_24!==16'h0011) $display("ERROR! at (9,24)\n");
if(pixels_10_24!==16'hff86) $display("ERROR! at (10,24)\n");
if(pixels_11_24!==16'hfe88) $display("ERROR! at (11,24)\n");
if(pixels_12_24!==16'hfd38) $display("ERROR! at (12,24)\n");
if(pixels_13_24!==16'hfe21) $display("ERROR! at (13,24)\n");
if(pixels_14_24!==16'hff8a) $display("ERROR! at (14,24)\n");
if(pixels_15_24!==16'h0567) $display("ERROR! at (15,24)\n");
if(pixels_16_24!==16'h0277) $display("ERROR! at (16,24)\n");
if(pixels_17_24!==16'h0091) $display("ERROR! at (17,24)\n");
if(pixels_18_24!==16'hf8e6) $display("ERROR! at (18,24)\n");
if(pixels_19_24!==16'hf5b4) $display("ERROR! at (19,24)\n");
if(pixels_20_24!==16'h015f) $display("ERROR! at (20,24)\n");
if(pixels_21_24!==16'hffac) $display("ERROR! at (21,24)\n");
if(pixels_22_24!==16'h0074) $display("ERROR! at (22,24)\n");
if(pixels_23_24!==16'hfcda) $display("ERROR! at (23,24)\n");
if(pixels_24_24!==16'hfb53) $display("ERROR! at (24,24)\n");
if(pixels_25_24!==16'h016b) $display("ERROR! at (25,24)\n");
if(pixels_26_24!==16'h038a) $display("ERROR! at (26,24)\n");
if(pixels_27_24!==16'h00bb) $display("ERROR! at (27,24)\n");
if(pixels_28_24!==16'hfc1e) $display("ERROR! at (28,24)\n");
if(pixels_29_24!==16'h02b4) $display("ERROR! at (29,24)\n");
if(pixels_30_24!==16'h0558) $display("ERROR! at (30,24)\n");
if(pixels_31_24!==16'hffd2) $display("ERROR! at (31,24)\n");
if(pixels_0_25!==16'hff82) $display("ERROR! at (0,25)\n");
if(pixels_1_25!==16'hfea3) $display("ERROR! at (1,25)\n");
if(pixels_2_25!==16'hfbab) $display("ERROR! at (2,25)\n");
if(pixels_3_25!==16'hfd56) $display("ERROR! at (3,25)\n");
if(pixels_4_25!==16'hfbbd) $display("ERROR! at (4,25)\n");
if(pixels_5_25!==16'h05be) $display("ERROR! at (5,25)\n");
if(pixels_6_25!==16'h07d3) $display("ERROR! at (6,25)\n");
if(pixels_7_25!==16'h066c) $display("ERROR! at (7,25)\n");
if(pixels_8_25!==16'h034c) $display("ERROR! at (8,25)\n");
if(pixels_9_25!==16'hfec7) $display("ERROR! at (9,25)\n");
if(pixels_10_25!==16'hfbf3) $display("ERROR! at (10,25)\n");
if(pixels_11_25!==16'hf733) $display("ERROR! at (11,25)\n");
if(pixels_12_25!==16'h02d1) $display("ERROR! at (12,25)\n");
if(pixels_13_25!==16'hfd30) $display("ERROR! at (13,25)\n");
if(pixels_14_25!==16'h0106) $display("ERROR! at (14,25)\n");
if(pixels_15_25!==16'hfac1) $display("ERROR! at (15,25)\n");
if(pixels_16_25!==16'hff6f) $display("ERROR! at (16,25)\n");
if(pixels_17_25!==16'hffe9) $display("ERROR! at (17,25)\n");
if(pixels_18_25!==16'hff64) $display("ERROR! at (18,25)\n");
if(pixels_19_25!==16'hf995) $display("ERROR! at (19,25)\n");
if(pixels_20_25!==16'hfcc0) $display("ERROR! at (20,25)\n");
if(pixels_21_25!==16'h06e5) $display("ERROR! at (21,25)\n");
if(pixels_22_25!==16'h0271) $display("ERROR! at (22,25)\n");
if(pixels_23_25!==16'h01a3) $display("ERROR! at (23,25)\n");
if(pixels_24_25!==16'hfb98) $display("ERROR! at (24,25)\n");
if(pixels_25_25!==16'hfd3c) $display("ERROR! at (25,25)\n");
if(pixels_26_25!==16'hfd73) $display("ERROR! at (26,25)\n");
if(pixels_27_25!==16'h0233) $display("ERROR! at (27,25)\n");
if(pixels_28_25!==16'h02e4) $display("ERROR! at (28,25)\n");
if(pixels_29_25!==16'h0057) $display("ERROR! at (29,25)\n");
if(pixels_30_25!==16'h0227) $display("ERROR! at (30,25)\n");
if(pixels_31_25!==16'hfe64) $display("ERROR! at (31,25)\n");
if(pixels_0_26!==16'h00f8) $display("ERROR! at (0,26)\n");
if(pixels_1_26!==16'h01bc) $display("ERROR! at (1,26)\n");
if(pixels_2_26!==16'h066b) $display("ERROR! at (2,26)\n");
if(pixels_3_26!==16'h0609) $display("ERROR! at (3,26)\n");
if(pixels_4_26!==16'h00bc) $display("ERROR! at (4,26)\n");
if(pixels_5_26!==16'hfeab) $display("ERROR! at (5,26)\n");
if(pixels_6_26!==16'h052a) $display("ERROR! at (6,26)\n");
if(pixels_7_26!==16'hfe70) $display("ERROR! at (7,26)\n");
if(pixels_8_26!==16'h0072) $display("ERROR! at (8,26)\n");
if(pixels_9_26!==16'hfc97) $display("ERROR! at (9,26)\n");
if(pixels_10_26!==16'h08f3) $display("ERROR! at (10,26)\n");
if(pixels_11_26!==16'h036e) $display("ERROR! at (11,26)\n");
if(pixels_12_26!==16'h006d) $display("ERROR! at (12,26)\n");
if(pixels_13_26!==16'h0076) $display("ERROR! at (13,26)\n");
if(pixels_14_26!==16'hfd9f) $display("ERROR! at (14,26)\n");
if(pixels_15_26!==16'h0277) $display("ERROR! at (15,26)\n");
if(pixels_16_26!==16'h044e) $display("ERROR! at (16,26)\n");
if(pixels_17_26!==16'hfc98) $display("ERROR! at (17,26)\n");
if(pixels_18_26!==16'hfe44) $display("ERROR! at (18,26)\n");
if(pixels_19_26!==16'hf953) $display("ERROR! at (19,26)\n");
if(pixels_20_26!==16'hf97a) $display("ERROR! at (20,26)\n");
if(pixels_21_26!==16'hfec7) $display("ERROR! at (21,26)\n");
if(pixels_22_26!==16'hfec3) $display("ERROR! at (22,26)\n");
if(pixels_23_26!==16'hfa17) $display("ERROR! at (23,26)\n");
if(pixels_24_26!==16'hfd8a) $display("ERROR! at (24,26)\n");
if(pixels_25_26!==16'h0288) $display("ERROR! at (25,26)\n");
if(pixels_26_26!==16'h0002) $display("ERROR! at (26,26)\n");
if(pixels_27_26!==16'h0373) $display("ERROR! at (27,26)\n");
if(pixels_28_26!==16'h0059) $display("ERROR! at (28,26)\n");
if(pixels_29_26!==16'h01f2) $display("ERROR! at (29,26)\n");
if(pixels_30_26!==16'h01cd) $display("ERROR! at (30,26)\n");
if(pixels_31_26!==16'h01a5) $display("ERROR! at (31,26)\n");
if(pixels_0_27!==16'hfc9b) $display("ERROR! at (0,27)\n");
if(pixels_1_27!==16'hfee3) $display("ERROR! at (1,27)\n");
if(pixels_2_27!==16'hf84d) $display("ERROR! at (2,27)\n");
if(pixels_3_27!==16'h026a) $display("ERROR! at (3,27)\n");
if(pixels_4_27!==16'h03e0) $display("ERROR! at (4,27)\n");
if(pixels_5_27!==16'h0464) $display("ERROR! at (5,27)\n");
if(pixels_6_27!==16'h045a) $display("ERROR! at (6,27)\n");
if(pixels_7_27!==16'h00e9) $display("ERROR! at (7,27)\n");
if(pixels_8_27!==16'h0127) $display("ERROR! at (8,27)\n");
if(pixels_9_27!==16'h0018) $display("ERROR! at (9,27)\n");
if(pixels_10_27!==16'hf705) $display("ERROR! at (10,27)\n");
if(pixels_11_27!==16'hfeb0) $display("ERROR! at (11,27)\n");
if(pixels_12_27!==16'hfee2) $display("ERROR! at (12,27)\n");
if(pixels_13_27!==16'h091c) $display("ERROR! at (13,27)\n");
if(pixels_14_27!==16'hff75) $display("ERROR! at (14,27)\n");
if(pixels_15_27!==16'hfed5) $display("ERROR! at (15,27)\n");
if(pixels_16_27!==16'h02a4) $display("ERROR! at (16,27)\n");
if(pixels_17_27!==16'hffc7) $display("ERROR! at (17,27)\n");
if(pixels_18_27!==16'hfb9a) $display("ERROR! at (18,27)\n");
if(pixels_19_27!==16'hfdcd) $display("ERROR! at (19,27)\n");
if(pixels_20_27!==16'hffa3) $display("ERROR! at (20,27)\n");
if(pixels_21_27!==16'h0258) $display("ERROR! at (21,27)\n");
if(pixels_22_27!==16'h0433) $display("ERROR! at (22,27)\n");
if(pixels_23_27!==16'hfaa0) $display("ERROR! at (23,27)\n");
if(pixels_24_27!==16'hfb3f) $display("ERROR! at (24,27)\n");
if(pixels_25_27!==16'h06d4) $display("ERROR! at (25,27)\n");
if(pixels_26_27!==16'hfec8) $display("ERROR! at (26,27)\n");
if(pixels_27_27!==16'hfe6e) $display("ERROR! at (27,27)\n");
if(pixels_28_27!==16'h04e7) $display("ERROR! at (28,27)\n");
if(pixels_29_27!==16'hfe7f) $display("ERROR! at (29,27)\n");
if(pixels_30_27!==16'hfee8) $display("ERROR! at (30,27)\n");
if(pixels_31_27!==16'h01e6) $display("ERROR! at (31,27)\n");
if(pixels_0_28!==16'h01d7) $display("ERROR! at (0,28)\n");
if(pixels_1_28!==16'h0111) $display("ERROR! at (1,28)\n");
if(pixels_2_28!==16'h0222) $display("ERROR! at (2,28)\n");
if(pixels_3_28!==16'hfdb2) $display("ERROR! at (3,28)\n");
if(pixels_4_28!==16'h053b) $display("ERROR! at (4,28)\n");
if(pixels_5_28!==16'hfab3) $display("ERROR! at (5,28)\n");
if(pixels_6_28!==16'hfbc0) $display("ERROR! at (6,28)\n");
if(pixels_7_28!==16'hfe0e) $display("ERROR! at (7,28)\n");
if(pixels_8_28!==16'hfd40) $display("ERROR! at (8,28)\n");
if(pixels_9_28!==16'h038e) $display("ERROR! at (9,28)\n");
if(pixels_10_28!==16'h0046) $display("ERROR! at (10,28)\n");
if(pixels_11_28!==16'h0271) $display("ERROR! at (11,28)\n");
if(pixels_12_28!==16'h02d3) $display("ERROR! at (12,28)\n");
if(pixels_13_28!==16'hfdb8) $display("ERROR! at (13,28)\n");
if(pixels_14_28!==16'hff70) $display("ERROR! at (14,28)\n");
if(pixels_15_28!==16'h00a2) $display("ERROR! at (15,28)\n");
if(pixels_16_28!==16'h0240) $display("ERROR! at (16,28)\n");
if(pixels_17_28!==16'h0357) $display("ERROR! at (17,28)\n");
if(pixels_18_28!==16'h008a) $display("ERROR! at (18,28)\n");
if(pixels_19_28!==16'hfd61) $display("ERROR! at (19,28)\n");
if(pixels_20_28!==16'h02ea) $display("ERROR! at (20,28)\n");
if(pixels_21_28!==16'hffba) $display("ERROR! at (21,28)\n");
if(pixels_22_28!==16'h0112) $display("ERROR! at (22,28)\n");
if(pixels_23_28!==16'h0228) $display("ERROR! at (23,28)\n");
if(pixels_24_28!==16'hfd68) $display("ERROR! at (24,28)\n");
if(pixels_25_28!==16'hfda8) $display("ERROR! at (25,28)\n");
if(pixels_26_28!==16'h0aa9) $display("ERROR! at (26,28)\n");
if(pixels_27_28!==16'h010a) $display("ERROR! at (27,28)\n");
if(pixels_28_28!==16'h01a9) $display("ERROR! at (28,28)\n");
if(pixels_29_28!==16'h0201) $display("ERROR! at (29,28)\n");
if(pixels_30_28!==16'h02d7) $display("ERROR! at (30,28)\n");
if(pixels_31_28!==16'h013a) $display("ERROR! at (31,28)\n");
if(pixels_0_29!==16'hfeb5) $display("ERROR! at (0,29)\n");
if(pixels_1_29!==16'hff3b) $display("ERROR! at (1,29)\n");
if(pixels_2_29!==16'hfcfe) $display("ERROR! at (2,29)\n");
if(pixels_3_29!==16'h00d6) $display("ERROR! at (3,29)\n");
if(pixels_4_29!==16'h0283) $display("ERROR! at (4,29)\n");
if(pixels_5_29!==16'h0386) $display("ERROR! at (5,29)\n");
if(pixels_6_29!==16'hfe5f) $display("ERROR! at (6,29)\n");
if(pixels_7_29!==16'hfe1e) $display("ERROR! at (7,29)\n");
if(pixels_8_29!==16'hfecc) $display("ERROR! at (8,29)\n");
if(pixels_9_29!==16'hfbcb) $display("ERROR! at (9,29)\n");
if(pixels_10_29!==16'h05b4) $display("ERROR! at (10,29)\n");
if(pixels_11_29!==16'hfd0b) $display("ERROR! at (11,29)\n");
if(pixels_12_29!==16'h03cc) $display("ERROR! at (12,29)\n");
if(pixels_13_29!==16'h0536) $display("ERROR! at (13,29)\n");
if(pixels_14_29!==16'h0605) $display("ERROR! at (14,29)\n");
if(pixels_15_29!==16'hff61) $display("ERROR! at (15,29)\n");
if(pixels_16_29!==16'hfbfd) $display("ERROR! at (16,29)\n");
if(pixels_17_29!==16'hffc2) $display("ERROR! at (17,29)\n");
if(pixels_18_29!==16'h0049) $display("ERROR! at (18,29)\n");
if(pixels_19_29!==16'hfa17) $display("ERROR! at (19,29)\n");
if(pixels_20_29!==16'h0142) $display("ERROR! at (20,29)\n");
if(pixels_21_29!==16'h038b) $display("ERROR! at (21,29)\n");
if(pixels_22_29!==16'h038d) $display("ERROR! at (22,29)\n");
if(pixels_23_29!==16'h00cd) $display("ERROR! at (23,29)\n");
if(pixels_24_29!==16'h0094) $display("ERROR! at (24,29)\n");
if(pixels_25_29!==16'h0250) $display("ERROR! at (25,29)\n");
if(pixels_26_29!==16'h0406) $display("ERROR! at (26,29)\n");
if(pixels_27_29!==16'h0261) $display("ERROR! at (27,29)\n");
if(pixels_28_29!==16'hf703) $display("ERROR! at (28,29)\n");
if(pixels_29_29!==16'h03d3) $display("ERROR! at (29,29)\n");
if(pixels_30_29!==16'h0213) $display("ERROR! at (30,29)\n");
if(pixels_31_29!==16'hffa3) $display("ERROR! at (31,29)\n");
if(pixels_0_30!==16'h017c) $display("ERROR! at (0,30)\n");
if(pixels_1_30!==16'h0229) $display("ERROR! at (1,30)\n");
if(pixels_2_30!==16'h0035) $display("ERROR! at (2,30)\n");
if(pixels_3_30!==16'hfe92) $display("ERROR! at (3,30)\n");
if(pixels_4_30!==16'hfe19) $display("ERROR! at (4,30)\n");
if(pixels_5_30!==16'hfe52) $display("ERROR! at (5,30)\n");
if(pixels_6_30!==16'hfbe3) $display("ERROR! at (6,30)\n");
if(pixels_7_30!==16'hfd90) $display("ERROR! at (7,30)\n");
if(pixels_8_30!==16'h026b) $display("ERROR! at (8,30)\n");
if(pixels_9_30!==16'h00da) $display("ERROR! at (9,30)\n");
if(pixels_10_30!==16'hfe7b) $display("ERROR! at (10,30)\n");
if(pixels_11_30!==16'hff20) $display("ERROR! at (11,30)\n");
if(pixels_12_30!==16'h0024) $display("ERROR! at (12,30)\n");
if(pixels_13_30!==16'h0035) $display("ERROR! at (13,30)\n");
if(pixels_14_30!==16'hff62) $display("ERROR! at (14,30)\n");
if(pixels_15_30!==16'h019c) $display("ERROR! at (15,30)\n");
if(pixels_16_30!==16'h01a1) $display("ERROR! at (16,30)\n");
if(pixels_17_30!==16'h004f) $display("ERROR! at (17,30)\n");
if(pixels_18_30!==16'hffd6) $display("ERROR! at (18,30)\n");
if(pixels_19_30!==16'h009e) $display("ERROR! at (19,30)\n");
if(pixels_20_30!==16'h0028) $display("ERROR! at (20,30)\n");
if(pixels_21_30!==16'hffd6) $display("ERROR! at (21,30)\n");
if(pixels_22_30!==16'hff73) $display("ERROR! at (22,30)\n");
if(pixels_23_30!==16'hff13) $display("ERROR! at (23,30)\n");
if(pixels_24_30!==16'h0394) $display("ERROR! at (24,30)\n");
if(pixels_25_30!==16'hfeff) $display("ERROR! at (25,30)\n");
if(pixels_26_30!==16'h023a) $display("ERROR! at (26,30)\n");
if(pixels_27_30!==16'h05b2) $display("ERROR! at (27,30)\n");
if(pixels_28_30!==16'h05c9) $display("ERROR! at (28,30)\n");
if(pixels_29_30!==16'hff22) $display("ERROR! at (29,30)\n");
if(pixels_30_30!==16'h01d6) $display("ERROR! at (30,30)\n");
if(pixels_31_30!==16'h00ab) $display("ERROR! at (31,30)\n");
if(pixels_0_31!==16'h0000) $display("ERROR! at (0,31)\n");
if(pixels_1_31!==16'hff74) $display("ERROR! at (1,31)\n");
if(pixels_2_31!==16'h00d2) $display("ERROR! at (2,31)\n");
if(pixels_3_31!==16'h01ca) $display("ERROR! at (3,31)\n");
if(pixels_4_31!==16'h03c7) $display("ERROR! at (4,31)\n");
if(pixels_5_31!==16'hff9f) $display("ERROR! at (5,31)\n");
if(pixels_6_31!==16'hfeee) $display("ERROR! at (6,31)\n");
if(pixels_7_31!==16'hfde8) $display("ERROR! at (7,31)\n");
if(pixels_8_31!==16'hff74) $display("ERROR! at (8,31)\n");
if(pixels_9_31!==16'h00df) $display("ERROR! at (9,31)\n");
if(pixels_10_31!==16'h0087) $display("ERROR! at (10,31)\n");
if(pixels_11_31!==16'h034e) $display("ERROR! at (11,31)\n");
if(pixels_12_31!==16'h013f) $display("ERROR! at (12,31)\n");
if(pixels_13_31!==16'h023e) $display("ERROR! at (13,31)\n");
if(pixels_14_31!==16'h00c4) $display("ERROR! at (14,31)\n");
if(pixels_15_31!==16'hfe75) $display("ERROR! at (15,31)\n");
if(pixels_16_31!==16'hfd9b) $display("ERROR! at (16,31)\n");
if(pixels_17_31!==16'hfefa) $display("ERROR! at (17,31)\n");
if(pixels_18_31!==16'hff55) $display("ERROR! at (18,31)\n");
if(pixels_19_31!==16'hff27) $display("ERROR! at (19,31)\n");
if(pixels_20_31!==16'hfed5) $display("ERROR! at (20,31)\n");
if(pixels_21_31!==16'h00bd) $display("ERROR! at (21,31)\n");
if(pixels_22_31!==16'h0162) $display("ERROR! at (22,31)\n");
if(pixels_23_31!==16'h007e) $display("ERROR! at (23,31)\n");
if(pixels_24_31!==16'h002a) $display("ERROR! at (24,31)\n");
if(pixels_25_31!==16'hff85) $display("ERROR! at (25,31)\n");
if(pixels_26_31!==16'h0251) $display("ERROR! at (26,31)\n");
if(pixels_27_31!==16'hfdb8) $display("ERROR! at (27,31)\n");
if(pixels_28_31!==16'hfebd) $display("ERROR! at (28,31)\n");
if(pixels_29_31!==16'hfdc5) $display("ERROR! at (29,31)\n");
if(pixels_30_31!==16'h048b) $display("ERROR! at (30,31)\n");
if(pixels_31_31!==16'h0190) $display("ERROR! at (31,31)\n");

    $finish;
    
end




always #5 clk = ~clk;

conv #(
    .col_length(col_length), 
    .word_length(word_length), 
    .double_word_length(double_word_length), 
    .kernel_size(kernel_size), 
    .image_size(image_size)
) u1 (
    .clk(clk),
    .rst(rst),
    .in_valid(in_valid),
    .weight_value(weight_value),
    .data_in(data_in),
    .data_out(data_out),
    .out_valid()
);

endmodule
