`timescale 1ns/1ns
module PE_tb_28();


parameter col_length = 8;
parameter word_length = 8;
parameter double_word_length = 16;
parameter kernel_size = 5;
parameter image_size = 28;


reg clk,rst,in_valid;

wire out_valid;
//weight in
reg [6272-1 :0] pe_input_feature_value='h04_09_f1_23_fe_fc_f8_03_fe_1a_17_07_0e_1d_05_f9_1e_f6_fd_fb_01_02_13_0e_05_11_ee_09_f7_fb_14_1d_ff_0f_ec_e4_eb_ed_f7_ef_19_dc_05_00_16_fb_ff_fe_04_f3_05_ef_f7_0d_04_02_fe_08_0a_ee_12_ef_ff_fb_11_fc_ff_03_e3_11_11_08_09_09_f6_07_f9_ef_00_ef_0a_0b_1a_07_0e_1a_00_f0_01_f5_07_00_ed_f1_f1_f8_0e_07_01_02_0f_d2_fe_0b_01_08_07_f3_fb_ee_e6_05_13_02_f3_0b_0a_04_09_0f_05_0c_f7_e3_f3_fa_f1_fe_0c_f2_11_ea_e2_f5_05_09_0d_06_f8_ef_f0_00_0c_e4_21_02_18_e5_19_08_fa_f2_0a_08_07_ef_04_04_02_0f_f3_f8_f3_f1_e7_f3_1d_0c_fb_e8_f5_ff_f6_00_0c_fa_e6_e3_fb_f7_fd_f7_e7_f9_f8_05_13_ee_09_f0_07_01_03_f5_11_f5_21_21_e3_e4_00_00_06_ed_ef_02_fc_f9_0d_fc_ff_07_08_f7_03_f3_fa_f8_fc_07_eb_f6_0b_ef_0d_0a_20_ed_fd_fd_0b_1e_00_fd_07_ff_eb_03_24_ff_f7_11_05_18_f8_e6_1f_05_0b_f0_ee_ed_04_17_f5_e5_03_04_0c_0a_fd_f6_ff_d2_f3_07_05_fd_01_e7_f5_f7_f9_15_f2_08_02_03_f9_15_0a_0f_06_04_25_0c_fe_0a_ff_e0_07_e9_07_09_0e_04_0e_08_0b_14_0b_f2_fd_0e_0a_f3_0e_ef_da_fb_f4_04_fc_f1_0a_11_0c_1d_20_fc_07_04_fb_0b_1f_15_09_f1_00_fa_16_f3_00_08_01_13_06_f9_09_fa_02_16_f0_0f_ff_fe_f5_02_29_f6_ec_f9_0a_e9_e3_10_2b_fd_02_f7_09_28_24_0b_f8_04_19_f2_f1_0f_e9_0d_df_f7_f2_f8_ff_eb_0f_03_fc_05_fe_e4_02_f4_f1_ed_f3_16_f6_01_f2_f6_02_06_fc_03_f9_fe_e7_06_1f_0b_05_14_1e_00_00_fb_eb_fc_fa_e0_0f_f6_de_0c_07_02_fc_ff_f2_0f_04_f8_f9_04_27_0f_06_18_f9_f6_06_ea_0d_02_0a_18_06_f3_fc_0f_0d_f2_0d_10_0c_0b_06_f0_0b_d6_12_f3_12_19_13_e5_f1_0d_0f_fa_0b_e8_eb_0c_04_1a_08_ea_ec_fe_03_ea_1f_10_f6_e9_1a_ff_05_fb_ea_23_26_f5_11_e5_fd_0d_05_f4_0b_04_f6_00_0e_f0_f7_fd_ee_1a_f8_10_0b_08_eb_0f_f5_15_0c_06_11_08_14_e8_1d_f3_f2_fa_f9_02_fd_11_0b_e7_f8_fc_e2_fd_16_04_1b_e9_15_00_fa_fc_03_08_0d_f8_05_0a_f1_f5_f2_02_f5_01_00_08_f7_02_27_06_ff_07_fa_f8_fa_05_15_00_0a_fc_ed_1b_20_2c_08_e8_f1_05_14_10_fa_14_f8_fb_fe_18_f9_10_10_e3_e7_07_01_00_03_00_fd_fa_06_01_03_15_fd_eb_f1_04_08_f5_1b_f1_15_00_04_f5_d8_f3_0e_fb_02_0d_0d_1b_f0_05_e6_07_04_17_f3_ef_37_10_ff_fb_0d_f9_f7_05_11_0f_0c_06_1c_04_01_ed_c8_f6_1b_01_17_02_fc_1f_1b_14_07_13_03_06_00_fa_f0_13_f3_08_0a_1f_f6_0e_fd_04_f0_00_10_06_f7_0c_17_05_f4_00_02_ff_f4_04_e8_d3_ff_e0_02_fe_f1_e8_f2_00_04_e3_01_09_0c_0b_e0_fe_1f_1a_f6_07_ed_fa_f1_fe_e9_fa_19_fe_0d_f1_0b_f3_fd_eb_1d_e0_fe_e2_1d_13_02_e8_03_f8_ff_f6_f1_ee_ea_f3_fc_10_fe_ed_15_fe_fe_e4_f5_ff_fa_0e_e2_03_e4_e0_0a_f3_10_f6_0a_fd_f3_f7_17_05_fc_0c_06_04_fc_02_f6_fd_0a_e2_07_0e_21_0c_11_ea_10_11_00_f7_ed_fe;
reg [224-1 :0] pe_input_weight_value='h00_00_00_25_0e_0b_ef_0f_29_e6_de_04_f3_03_f7_10_ef_f6_fb_05_15_16_01_f8_00_0a_00_ee;
reg [6272-1 :0] pe_input_feature_cols='b00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000_00011011_00011010_00011001_00011000_00010111_00010110_00010101_00010100_00010011_00010010_00010001_00010000_00001111_00001110_00001101_00001100_00001011_00001010_00001001_00001000_00000111_00000110_00000101_00000100_00000011_00000010_00000001_00000000;
reg [6272-1 :0] pe_input_feature_rows='b00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011011_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011010_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011001_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010111_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010110_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010101_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010100_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010011_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010010_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010001_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00010000_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001111_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001110_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001101_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001011_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001010_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001001_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000111_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000110_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000100_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000011_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000010_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
reg [224-1 :0] pe_input_weight_cols='b00000000_00000000_00000000_00000100_00000011_00000010_00000001_00000000_00000100_00000011_00000010_00000001_00000000_00000100_00000011_00000010_00000001_00000000_00000100_00000011_00000010_00000001_00000000_00000100_00000011_00000010_00000001_00000000;
reg [224-1 :0] pe_input_weight_rows='b00000000_00000000_00000000_00000100_00000100_00000100_00000100_00000100_00000011_00000011_00000011_00000011_00000011_00000010_00000010_00000010_00000010_00000010_00000001_00000001_00000001_00000001_00000001_00000000_00000000_00000000_00000000_00000000;

//pixel data
reg [double_word_length-1:0] feature_valid_num,weight_valid_num;

//for test only
reg [32*32*word_length*2-1:0] result;
wire signed [word_length*2*16 -1:0]data_out;
wire signed [col_length*16 -1:0]data_out_cols;
wire signed [col_length*16 -1:0]data_out_rows;

wire signed [word_length*2-1:0] answer_1_1,answer_1_2,answer_1_3,answer_1_4,answer_2_1,answer_2_2,answer_2_3,answer_2_4;
wire signed [word_length*2-1:0] answer_3_1,answer_3_2,answer_3_3,answer_3_4,answer_4_1,answer_4_2,answer_4_3,answer_4_4; 
wire signed [col_length-1:0] col_answer_1_1,col_answer_1_2,col_answer_1_3,col_answer_1_4,col_answer_2_1,col_answer_2_2,col_answer_2_3,col_answer_2_4,col_answer_3_1,col_answer_3_2,col_answer_3_3,col_answer_3_4,col_answer_4_1,col_answer_4_2,col_answer_4_3,col_answer_4_4; 
wire signed [col_length-1:0] row_answer_1_1,row_answer_1_2,row_answer_1_3,row_answer_1_4,row_answer_2_1,row_answer_2_2,row_answer_2_3,row_answer_2_4,row_answer_3_1,row_answer_3_2,row_answer_3_3,row_answer_3_4,row_answer_4_1,row_answer_4_2,row_answer_4_3,row_answer_4_4; 

assign {col_answer_4_4,col_answer_4_3,col_answer_4_2,col_answer_4_1, col_answer_3_4,col_answer_3_3,col_answer_3_2,col_answer_3_1, col_answer_2_4,col_answer_2_3,col_answer_2_2,col_answer_2_1, col_answer_1_4,col_answer_1_3,col_answer_1_2,col_answer_1_1}= data_out_cols;
assign {row_answer_4_4,row_answer_4_3,row_answer_4_2,row_answer_4_1, row_answer_3_4,row_answer_3_3,row_answer_3_2,row_answer_3_1, row_answer_2_4,row_answer_2_3,row_answer_2_2,row_answer_2_1, row_answer_1_4,row_answer_1_3,row_answer_1_2,row_answer_1_1}= data_out_rows;

assign {{answer_1_4},{answer_1_3},{answer_1_2},{answer_1_1}} = data_out[word_length*2*4 -1 -:word_length*2*4];
assign {{answer_2_4},{answer_2_3},{answer_2_2},{answer_2_1}} = data_out[word_length*2*8 -1 -:word_length*2*4];
assign {{answer_3_4},{answer_3_3},{answer_3_2},{answer_3_1}} = data_out[word_length*2*12 -1 -:word_length*2*4];
assign {{answer_4_4},{answer_4_3},{answer_4_2},{answer_4_1}} = data_out[word_length*2*16 -1 -:word_length*2*4];

wire signed  [word_length*2-1:0] pixels_0_0, pixels_0_1, pixels_0_2, pixels_0_3, pixels_0_4, pixels_0_5, pixels_0_6, pixels_0_7, pixels_0_8, pixels_0_9, pixels_0_10, pixels_0_11, pixels_0_12, pixels_0_13, pixels_0_14, pixels_0_15, pixels_0_16, pixels_0_17, pixels_0_18, pixels_0_19, pixels_0_20, pixels_0_21, pixels_0_22, pixels_0_23, pixels_0_24, pixels_0_25, pixels_0_26, pixels_0_27, pixels_0_28, pixels_0_29, pixels_0_30, pixels_0_31, pixels_1_0, pixels_1_1, pixels_1_2, pixels_1_3, pixels_1_4, pixels_1_5, pixels_1_6, pixels_1_7, pixels_1_8, pixels_1_9, pixels_1_10, pixels_1_11, pixels_1_12, pixels_1_13, pixels_1_14, pixels_1_15, pixels_1_16, pixels_1_17, pixels_1_18, pixels_1_19, pixels_1_20, pixels_1_21, pixels_1_22, pixels_1_23, pixels_1_24, pixels_1_25, pixels_1_26, pixels_1_27, pixels_1_28, pixels_1_29, pixels_1_30, pixels_1_31, pixels_2_0, pixels_2_1, pixels_2_2, pixels_2_3, pixels_2_4, pixels_2_5, pixels_2_6, pixels_2_7, pixels_2_8, pixels_2_9, pixels_2_10, pixels_2_11, pixels_2_12, pixels_2_13, pixels_2_14, pixels_2_15, pixels_2_16, pixels_2_17, pixels_2_18, pixels_2_19, pixels_2_20, pixels_2_21, pixels_2_22, pixels_2_23, pixels_2_24, pixels_2_25, pixels_2_26, pixels_2_27, pixels_2_28, pixels_2_29, pixels_2_30, pixels_2_31, pixels_3_0, pixels_3_1, pixels_3_2, pixels_3_3, pixels_3_4, pixels_3_5, pixels_3_6, pixels_3_7, pixels_3_8, pixels_3_9, pixels_3_10, pixels_3_11, pixels_3_12, pixels_3_13, pixels_3_14, pixels_3_15, pixels_3_16, pixels_3_17, pixels_3_18, pixels_3_19, pixels_3_20, pixels_3_21, pixels_3_22, pixels_3_23, pixels_3_24, pixels_3_25, pixels_3_26, pixels_3_27, pixels_3_28, pixels_3_29, pixels_3_30, pixels_3_31, pixels_4_0, pixels_4_1, pixels_4_2, pixels_4_3, pixels_4_4, pixels_4_5, pixels_4_6, pixels_4_7, pixels_4_8, pixels_4_9, pixels_4_10, pixels_4_11, pixels_4_12, pixels_4_13, pixels_4_14, pixels_4_15, pixels_4_16, pixels_4_17, pixels_4_18, pixels_4_19, pixels_4_20, pixels_4_21, pixels_4_22, pixels_4_23, pixels_4_24, pixels_4_25, pixels_4_26, pixels_4_27, pixels_4_28, pixels_4_29, pixels_4_30, pixels_4_31, pixels_5_0, pixels_5_1, pixels_5_2, pixels_5_3, pixels_5_4, pixels_5_5, pixels_5_6, pixels_5_7, pixels_5_8, pixels_5_9, pixels_5_10, pixels_5_11, pixels_5_12, pixels_5_13, pixels_5_14, pixels_5_15, pixels_5_16, pixels_5_17, pixels_5_18, pixels_5_19, pixels_5_20, pixels_5_21, pixels_5_22, pixels_5_23, pixels_5_24, pixels_5_25, pixels_5_26, pixels_5_27, pixels_5_28, pixels_5_29, pixels_5_30, pixels_5_31, pixels_6_0, pixels_6_1, pixels_6_2, pixels_6_3, pixels_6_4, pixels_6_5, pixels_6_6, pixels_6_7, pixels_6_8, pixels_6_9, pixels_6_10, pixels_6_11, pixels_6_12, pixels_6_13, pixels_6_14, pixels_6_15, pixels_6_16, pixels_6_17, pixels_6_18, pixels_6_19, pixels_6_20, pixels_6_21, pixels_6_22, pixels_6_23, pixels_6_24, pixels_6_25, pixels_6_26, pixels_6_27, pixels_6_28, pixels_6_29, pixels_6_30, pixels_6_31, pixels_7_0, pixels_7_1, pixels_7_2, pixels_7_3, pixels_7_4, pixels_7_5, pixels_7_6, pixels_7_7, pixels_7_8, pixels_7_9, pixels_7_10, pixels_7_11, pixels_7_12, pixels_7_13, pixels_7_14, pixels_7_15, pixels_7_16, pixels_7_17, pixels_7_18, pixels_7_19, pixels_7_20, pixels_7_21, pixels_7_22, pixels_7_23, pixels_7_24, pixels_7_25, pixels_7_26, pixels_7_27, pixels_7_28, pixels_7_29, pixels_7_30, pixels_7_31, pixels_8_0, pixels_8_1, pixels_8_2, pixels_8_3, pixels_8_4, pixels_8_5, pixels_8_6, pixels_8_7, pixels_8_8, pixels_8_9, pixels_8_10, pixels_8_11, pixels_8_12, pixels_8_13, pixels_8_14, pixels_8_15, pixels_8_16, pixels_8_17, pixels_8_18, pixels_8_19, pixels_8_20, pixels_8_21, pixels_8_22, pixels_8_23, pixels_8_24, pixels_8_25, pixels_8_26, pixels_8_27, pixels_8_28, pixels_8_29, pixels_8_30, pixels_8_31, pixels_9_0, pixels_9_1, pixels_9_2, pixels_9_3, pixels_9_4, pixels_9_5, pixels_9_6, pixels_9_7, pixels_9_8, pixels_9_9, pixels_9_10, pixels_9_11, pixels_9_12, pixels_9_13, pixels_9_14, pixels_9_15, pixels_9_16, pixels_9_17, pixels_9_18, pixels_9_19, pixels_9_20, pixels_9_21, pixels_9_22, pixels_9_23, pixels_9_24, pixels_9_25, pixels_9_26, pixels_9_27, pixels_9_28, pixels_9_29, pixels_9_30, pixels_9_31, pixels_10_0, pixels_10_1, pixels_10_2, pixels_10_3, pixels_10_4, pixels_10_5, pixels_10_6, pixels_10_7, pixels_10_8, pixels_10_9, pixels_10_10, pixels_10_11, pixels_10_12, pixels_10_13, pixels_10_14, pixels_10_15, pixels_10_16, pixels_10_17, pixels_10_18, pixels_10_19, pixels_10_20, pixels_10_21, pixels_10_22, pixels_10_23, pixels_10_24, pixels_10_25, pixels_10_26, pixels_10_27, pixels_10_28, pixels_10_29, pixels_10_30, pixels_10_31, pixels_11_0, pixels_11_1, pixels_11_2, pixels_11_3, pixels_11_4, pixels_11_5, pixels_11_6, pixels_11_7, pixels_11_8, pixels_11_9, pixels_11_10, pixels_11_11, pixels_11_12, pixels_11_13, pixels_11_14, pixels_11_15, pixels_11_16, pixels_11_17, pixels_11_18, pixels_11_19, pixels_11_20, pixels_11_21, pixels_11_22, pixels_11_23, pixels_11_24, pixels_11_25, pixels_11_26, pixels_11_27, pixels_11_28, pixels_11_29, pixels_11_30, pixels_11_31, pixels_12_0, pixels_12_1, pixels_12_2, pixels_12_3, pixels_12_4, pixels_12_5, pixels_12_6, pixels_12_7, pixels_12_8, pixels_12_9, pixels_12_10, pixels_12_11, pixels_12_12, pixels_12_13, pixels_12_14, pixels_12_15, pixels_12_16, pixels_12_17, pixels_12_18, pixels_12_19, pixels_12_20, pixels_12_21, pixels_12_22, pixels_12_23, pixels_12_24, pixels_12_25, pixels_12_26, pixels_12_27, pixels_12_28, pixels_12_29, pixels_12_30, pixels_12_31, pixels_13_0, pixels_13_1, pixels_13_2, pixels_13_3, pixels_13_4, pixels_13_5, pixels_13_6, pixels_13_7, pixels_13_8, pixels_13_9, pixels_13_10, pixels_13_11, pixels_13_12, pixels_13_13, pixels_13_14, pixels_13_15, pixels_13_16, pixels_13_17, pixels_13_18, pixels_13_19, pixels_13_20, pixels_13_21, pixels_13_22, pixels_13_23, pixels_13_24, pixels_13_25, pixels_13_26, pixels_13_27, pixels_13_28, pixels_13_29, pixels_13_30, pixels_13_31, pixels_14_0, pixels_14_1, pixels_14_2, pixels_14_3, pixels_14_4, pixels_14_5, pixels_14_6, pixels_14_7, pixels_14_8, pixels_14_9, pixels_14_10, pixels_14_11, pixels_14_12, pixels_14_13, pixels_14_14, pixels_14_15, pixels_14_16, pixels_14_17, pixels_14_18, pixels_14_19, pixels_14_20, pixels_14_21, pixels_14_22, pixels_14_23, pixels_14_24, pixels_14_25, pixels_14_26, pixels_14_27, pixels_14_28, pixels_14_29, pixels_14_30, pixels_14_31, pixels_15_0, pixels_15_1, pixels_15_2, pixels_15_3, pixels_15_4, pixels_15_5, pixels_15_6, pixels_15_7, pixels_15_8, pixels_15_9, pixels_15_10, pixels_15_11, pixels_15_12, pixels_15_13, pixels_15_14, pixels_15_15, pixels_15_16, pixels_15_17, pixels_15_18, pixels_15_19, pixels_15_20, pixels_15_21, pixels_15_22, pixels_15_23, pixels_15_24, pixels_15_25, pixels_15_26, pixels_15_27, pixels_15_28, pixels_15_29, pixels_15_30, pixels_15_31, pixels_16_0, pixels_16_1, pixels_16_2, pixels_16_3, pixels_16_4, pixels_16_5, pixels_16_6, pixels_16_7, pixels_16_8, pixels_16_9, pixels_16_10, pixels_16_11, pixels_16_12, pixels_16_13, pixels_16_14, pixels_16_15, pixels_16_16, pixels_16_17, pixels_16_18, pixels_16_19, pixels_16_20, pixels_16_21, pixels_16_22, pixels_16_23, pixels_16_24, pixels_16_25, pixels_16_26, pixels_16_27, pixels_16_28, pixels_16_29, pixels_16_30, pixels_16_31, pixels_17_0, pixels_17_1, pixels_17_2, pixels_17_3, pixels_17_4, pixels_17_5, pixels_17_6, pixels_17_7, pixels_17_8, pixels_17_9, pixels_17_10, pixels_17_11, pixels_17_12, pixels_17_13, pixels_17_14, pixels_17_15, pixels_17_16, pixels_17_17, pixels_17_18, pixels_17_19, pixels_17_20, pixels_17_21, pixels_17_22, pixels_17_23, pixels_17_24, pixels_17_25, pixels_17_26, pixels_17_27, pixels_17_28, pixels_17_29, pixels_17_30, pixels_17_31, pixels_18_0, pixels_18_1, pixels_18_2, pixels_18_3, pixels_18_4, pixels_18_5, pixels_18_6, pixels_18_7, pixels_18_8, pixels_18_9, pixels_18_10, pixels_18_11, pixels_18_12, pixels_18_13, pixels_18_14, pixels_18_15, pixels_18_16, pixels_18_17, pixels_18_18, pixels_18_19, pixels_18_20, pixels_18_21, pixels_18_22, pixels_18_23, pixels_18_24, pixels_18_25, pixels_18_26, pixels_18_27, pixels_18_28, pixels_18_29, pixels_18_30, pixels_18_31, pixels_19_0, pixels_19_1, pixels_19_2, pixels_19_3, pixels_19_4, pixels_19_5, pixels_19_6, pixels_19_7, pixels_19_8, pixels_19_9, pixels_19_10, pixels_19_11, pixels_19_12, pixels_19_13, pixels_19_14, pixels_19_15, pixels_19_16, pixels_19_17, pixels_19_18, pixels_19_19, pixels_19_20, pixels_19_21, pixels_19_22, pixels_19_23, pixels_19_24, pixels_19_25, pixels_19_26, pixels_19_27, pixels_19_28, pixels_19_29, pixels_19_30, pixels_19_31, pixels_20_0, pixels_20_1, pixels_20_2, pixels_20_3, pixels_20_4, pixels_20_5, pixels_20_6, pixels_20_7, pixels_20_8, pixels_20_9, pixels_20_10, pixels_20_11, pixels_20_12, pixels_20_13, pixels_20_14, pixels_20_15, pixels_20_16, pixels_20_17, pixels_20_18, pixels_20_19, pixels_20_20, pixels_20_21, pixels_20_22, pixels_20_23, pixels_20_24, pixels_20_25, pixels_20_26, pixels_20_27, pixels_20_28, pixels_20_29, pixels_20_30, pixels_20_31, pixels_21_0, pixels_21_1, pixels_21_2, pixels_21_3, pixels_21_4, pixels_21_5, pixels_21_6, pixels_21_7, pixels_21_8, pixels_21_9, pixels_21_10, pixels_21_11, pixels_21_12, pixels_21_13, pixels_21_14, pixels_21_15, pixels_21_16, pixels_21_17, pixels_21_18, pixels_21_19, pixels_21_20, pixels_21_21, pixels_21_22, pixels_21_23, pixels_21_24, pixels_21_25, pixels_21_26, pixels_21_27, pixels_21_28, pixels_21_29, pixels_21_30, pixels_21_31, pixels_22_0, pixels_22_1, pixels_22_2, pixels_22_3, pixels_22_4, pixels_22_5, pixels_22_6, pixels_22_7, pixels_22_8, pixels_22_9, pixels_22_10, pixels_22_11, pixels_22_12, pixels_22_13, pixels_22_14, pixels_22_15, pixels_22_16, pixels_22_17, pixels_22_18, pixels_22_19, pixels_22_20, pixels_22_21, pixels_22_22, pixels_22_23, pixels_22_24, pixels_22_25, pixels_22_26, pixels_22_27, pixels_22_28, pixels_22_29, pixels_22_30, pixels_22_31, 
pixels_23_0, pixels_23_1, pixels_23_2, pixels_23_3, pixels_23_4, pixels_23_5, pixels_23_6, pixels_23_7, pixels_23_8, pixels_23_9, pixels_23_10, pixels_23_11, pixels_23_12, pixels_23_13, pixels_23_14, pixels_23_15, pixels_23_16, pixels_23_17, pixels_23_18, pixels_23_19, pixels_23_20, pixels_23_21, pixels_23_22, pixels_23_23, pixels_23_24, pixels_23_25, pixels_23_26, pixels_23_27, pixels_23_28, pixels_23_29, pixels_23_30, pixels_23_31, pixels_24_0, pixels_24_1, pixels_24_2, pixels_24_3, pixels_24_4, pixels_24_5, pixels_24_6, pixels_24_7, pixels_24_8, pixels_24_9, pixels_24_10, pixels_24_11, pixels_24_12, pixels_24_13, pixels_24_14, pixels_24_15, pixels_24_16, pixels_24_17, pixels_24_18, pixels_24_19, pixels_24_20, pixels_24_21, pixels_24_22, pixels_24_23, pixels_24_24, pixels_24_25, pixels_24_26, pixels_24_27, pixels_24_28, pixels_24_29, pixels_24_30, pixels_24_31, pixels_25_0, pixels_25_1, pixels_25_2, pixels_25_3, pixels_25_4, pixels_25_5, pixels_25_6, pixels_25_7, pixels_25_8, pixels_25_9, pixels_25_10, pixels_25_11, pixels_25_12, pixels_25_13, pixels_25_14, pixels_25_15, pixels_25_16, pixels_25_17, pixels_25_18, pixels_25_19, pixels_25_20, pixels_25_21, pixels_25_22, pixels_25_23, pixels_25_24, pixels_25_25, pixels_25_26, pixels_25_27, pixels_25_28, pixels_25_29, pixels_25_30, pixels_25_31, pixels_26_0, pixels_26_1, pixels_26_2, pixels_26_3, pixels_26_4, pixels_26_5, pixels_26_6, pixels_26_7, pixels_26_8, pixels_26_9, pixels_26_10, pixels_26_11, pixels_26_12, pixels_26_13, pixels_26_14, pixels_26_15, pixels_26_16, pixels_26_17, pixels_26_18, pixels_26_19, pixels_26_20, pixels_26_21, pixels_26_22, pixels_26_23, pixels_26_24, pixels_26_25, pixels_26_26, pixels_26_27, pixels_26_28, pixels_26_29, pixels_26_30, pixels_26_31, pixels_27_0, pixels_27_1, pixels_27_2, pixels_27_3, pixels_27_4, pixels_27_5, pixels_27_6, pixels_27_7, pixels_27_8, pixels_27_9, pixels_27_10, pixels_27_11, pixels_27_12, pixels_27_13, pixels_27_14, pixels_27_15, pixels_27_16, pixels_27_17, pixels_27_18, pixels_27_19, pixels_27_20, pixels_27_21, pixels_27_22, pixels_27_23, pixels_27_24, pixels_27_25, pixels_27_26, pixels_27_27, pixels_27_28, pixels_27_29, pixels_27_30, pixels_27_31, pixels_28_0, pixels_28_1, pixels_28_2, pixels_28_3, pixels_28_4, pixels_28_5, pixels_28_6, pixels_28_7, pixels_28_8, pixels_28_9, pixels_28_10, pixels_28_11, pixels_28_12, pixels_28_13, pixels_28_14, pixels_28_15, pixels_28_16, pixels_28_17, pixels_28_18, pixels_28_19, pixels_28_20, pixels_28_21, pixels_28_22, pixels_28_23, pixels_28_24, pixels_28_25, pixels_28_26, pixels_28_27, pixels_28_28, pixels_28_29, pixels_28_30, pixels_28_31, pixels_29_0, pixels_29_1, pixels_29_2, pixels_29_3, pixels_29_4, pixels_29_5, pixels_29_6, pixels_29_7, pixels_29_8, pixels_29_9, pixels_29_10, pixels_29_11, pixels_29_12, pixels_29_13, pixels_29_14, pixels_29_15, pixels_29_16, pixels_29_17, pixels_29_18, pixels_29_19, pixels_29_20, pixels_29_21, pixels_29_22, pixels_29_23, pixels_29_24, pixels_29_25, pixels_29_26, pixels_29_27, pixels_29_28, pixels_29_29, pixels_29_30, pixels_29_31, pixels_30_0, pixels_30_1, pixels_30_2, pixels_30_3, pixels_30_4, pixels_30_5, pixels_30_6, pixels_30_7, pixels_30_8, pixels_30_9, pixels_30_10, pixels_30_11, pixels_30_12, pixels_30_13, pixels_30_14, pixels_30_15, pixels_30_16, pixels_30_17, pixels_30_18, pixels_30_19, pixels_30_20, pixels_30_21, pixels_30_22, pixels_30_23, pixels_30_24, pixels_30_25, pixels_30_26, pixels_30_27, pixels_30_28, pixels_30_29, pixels_30_30, pixels_30_31, pixels_31_0, pixels_31_1, pixels_31_2, pixels_31_3, pixels_31_4, pixels_31_5, pixels_31_6, pixels_31_7, pixels_31_8, pixels_31_9, pixels_31_10, pixels_31_11, pixels_31_12, pixels_31_13, pixels_31_14, pixels_31_15, pixels_31_16, pixels_31_17, pixels_31_18, pixels_31_19, pixels_31_20, pixels_31_21, pixels_31_22, pixels_31_23, pixels_31_24, pixels_31_25, pixels_31_26, pixels_31_27, pixels_31_28, pixels_31_29, pixels_31_30, pixels_31_31;

assign pixels_0_0 = {result[1*word_length*2-1 -: word_length*2]};
assign pixels_1_0 = {result[2*word_length*2-1 -: word_length*2]};
assign pixels_2_0 = {result[3*word_length*2-1 -: word_length*2]};
assign pixels_3_0 = {result[4*word_length*2-1 -: word_length*2]};
assign pixels_4_0 = {result[5*word_length*2-1 -: word_length*2]};
assign pixels_5_0 = {result[6*word_length*2-1 -: word_length*2]};
assign pixels_6_0 = {result[7*word_length*2-1 -: word_length*2]};
assign pixels_7_0 = {result[8*word_length*2-1 -: word_length*2]};
assign pixels_8_0 = {result[9*word_length*2-1 -: word_length*2]};
assign pixels_9_0 = {result[10*word_length*2-1 -: word_length*2]};
assign pixels_10_0 = {result[11*word_length*2-1 -: word_length*2]};
assign pixels_11_0 = {result[12*word_length*2-1 -: word_length*2]};
assign pixels_12_0 = {result[13*word_length*2-1 -: word_length*2]};
assign pixels_13_0 = {result[14*word_length*2-1 -: word_length*2]};
assign pixels_14_0 = {result[15*word_length*2-1 -: word_length*2]};
assign pixels_15_0 = {result[16*word_length*2-1 -: word_length*2]};
assign pixels_16_0 = {result[17*word_length*2-1 -: word_length*2]};
assign pixels_17_0 = {result[18*word_length*2-1 -: word_length*2]};
assign pixels_18_0 = {result[19*word_length*2-1 -: word_length*2]};
assign pixels_19_0 = {result[20*word_length*2-1 -: word_length*2]};
assign pixels_20_0 = {result[21*word_length*2-1 -: word_length*2]};
assign pixels_21_0 = {result[22*word_length*2-1 -: word_length*2]};
assign pixels_22_0 = {result[23*word_length*2-1 -: word_length*2]};
assign pixels_23_0 = {result[24*word_length*2-1 -: word_length*2]};
assign pixels_24_0 = {result[25*word_length*2-1 -: word_length*2]};
assign pixels_25_0 = {result[26*word_length*2-1 -: word_length*2]};
assign pixels_26_0 = {result[27*word_length*2-1 -: word_length*2]};
assign pixels_27_0 = {result[28*word_length*2-1 -: word_length*2]};
assign pixels_28_0 = {result[29*word_length*2-1 -: word_length*2]};
assign pixels_29_0 = {result[30*word_length*2-1 -: word_length*2]};
assign pixels_30_0 = {result[31*word_length*2-1 -: word_length*2]};
assign pixels_31_0 = {result[32*word_length*2-1 -: word_length*2]};
assign pixels_0_1 = {result[33*word_length*2-1 -: word_length*2]};
assign pixels_1_1 = {result[34*word_length*2-1 -: word_length*2]};
assign pixels_2_1 = {result[35*word_length*2-1 -: word_length*2]};
assign pixels_3_1 = {result[36*word_length*2-1 -: word_length*2]};
assign pixels_4_1 = {result[37*word_length*2-1 -: word_length*2]};
assign pixels_5_1 = {result[38*word_length*2-1 -: word_length*2]};
assign pixels_6_1 = {result[39*word_length*2-1 -: word_length*2]};
assign pixels_7_1 = {result[40*word_length*2-1 -: word_length*2]};
assign pixels_8_1 = {result[41*word_length*2-1 -: word_length*2]};
assign pixels_9_1 = {result[42*word_length*2-1 -: word_length*2]};
assign pixels_10_1 = {result[43*word_length*2-1 -: word_length*2]};
assign pixels_11_1 = {result[44*word_length*2-1 -: word_length*2]};
assign pixels_12_1 = {result[45*word_length*2-1 -: word_length*2]};
assign pixels_13_1 = {result[46*word_length*2-1 -: word_length*2]};
assign pixels_14_1 = {result[47*word_length*2-1 -: word_length*2]};
assign pixels_15_1 = {result[48*word_length*2-1 -: word_length*2]};
assign pixels_16_1 = {result[49*word_length*2-1 -: word_length*2]};
assign pixels_17_1 = {result[50*word_length*2-1 -: word_length*2]};
assign pixels_18_1 = {result[51*word_length*2-1 -: word_length*2]};
assign pixels_19_1 = {result[52*word_length*2-1 -: word_length*2]};
assign pixels_20_1 = {result[53*word_length*2-1 -: word_length*2]};
assign pixels_21_1 = {result[54*word_length*2-1 -: word_length*2]};
assign pixels_22_1 = {result[55*word_length*2-1 -: word_length*2]};
assign pixels_23_1 = {result[56*word_length*2-1 -: word_length*2]};
assign pixels_24_1 = {result[57*word_length*2-1 -: word_length*2]};
assign pixels_25_1 = {result[58*word_length*2-1 -: word_length*2]};
assign pixels_26_1 = {result[59*word_length*2-1 -: word_length*2]};
assign pixels_27_1 = {result[60*word_length*2-1 -: word_length*2]};
assign pixels_28_1 = {result[61*word_length*2-1 -: word_length*2]};
assign pixels_29_1 = {result[62*word_length*2-1 -: word_length*2]};
assign pixels_30_1 = {result[63*word_length*2-1 -: word_length*2]};
assign pixels_31_1 = {result[64*word_length*2-1 -: word_length*2]};
assign pixels_0_2 = {result[65*word_length*2-1 -: word_length*2]};
assign pixels_1_2 = {result[66*word_length*2-1 -: word_length*2]};
assign pixels_2_2 = {result[67*word_length*2-1 -: word_length*2]};
assign pixels_3_2 = {result[68*word_length*2-1 -: word_length*2]};
assign pixels_4_2 = {result[69*word_length*2-1 -: word_length*2]};
assign pixels_5_2 = {result[70*word_length*2-1 -: word_length*2]};
assign pixels_6_2 = {result[71*word_length*2-1 -: word_length*2]};
assign pixels_7_2 = {result[72*word_length*2-1 -: word_length*2]};
assign pixels_8_2 = {result[73*word_length*2-1 -: word_length*2]};
assign pixels_9_2 = {result[74*word_length*2-1 -: word_length*2]};
assign pixels_10_2 = {result[75*word_length*2-1 -: word_length*2]};
assign pixels_11_2 = {result[76*word_length*2-1 -: word_length*2]};
assign pixels_12_2 = {result[77*word_length*2-1 -: word_length*2]};
assign pixels_13_2 = {result[78*word_length*2-1 -: word_length*2]};
assign pixels_14_2 = {result[79*word_length*2-1 -: word_length*2]};
assign pixels_15_2 = {result[80*word_length*2-1 -: word_length*2]};
assign pixels_16_2 = {result[81*word_length*2-1 -: word_length*2]};
assign pixels_17_2 = {result[82*word_length*2-1 -: word_length*2]};
assign pixels_18_2 = {result[83*word_length*2-1 -: word_length*2]};
assign pixels_19_2 = {result[84*word_length*2-1 -: word_length*2]};
assign pixels_20_2 = {result[85*word_length*2-1 -: word_length*2]};
assign pixels_21_2 = {result[86*word_length*2-1 -: word_length*2]};
assign pixels_22_2 = {result[87*word_length*2-1 -: word_length*2]};
assign pixels_23_2 = {result[88*word_length*2-1 -: word_length*2]};
assign pixels_24_2 = {result[89*word_length*2-1 -: word_length*2]};
assign pixels_25_2 = {result[90*word_length*2-1 -: word_length*2]};
assign pixels_26_2 = {result[91*word_length*2-1 -: word_length*2]};
assign pixels_27_2 = {result[92*word_length*2-1 -: word_length*2]};
assign pixels_28_2 = {result[93*word_length*2-1 -: word_length*2]};
assign pixels_29_2 = {result[94*word_length*2-1 -: word_length*2]};
assign pixels_30_2 = {result[95*word_length*2-1 -: word_length*2]};
assign pixels_31_2 = {result[96*word_length*2-1 -: word_length*2]};
assign pixels_0_3 = {result[97*word_length*2-1 -: word_length*2]};
assign pixels_1_3 = {result[98*word_length*2-1 -: word_length*2]};
assign pixels_2_3 = {result[99*word_length*2-1 -: word_length*2]};
assign pixels_3_3 = {result[100*word_length*2-1 -: word_length*2]};
assign pixels_4_3 = {result[101*word_length*2-1 -: word_length*2]};
assign pixels_5_3 = {result[102*word_length*2-1 -: word_length*2]};
assign pixels_6_3 = {result[103*word_length*2-1 -: word_length*2]};
assign pixels_7_3 = {result[104*word_length*2-1 -: word_length*2]};
assign pixels_8_3 = {result[105*word_length*2-1 -: word_length*2]};
assign pixels_9_3 = {result[106*word_length*2-1 -: word_length*2]};
assign pixels_10_3 = {result[107*word_length*2-1 -: word_length*2]};
assign pixels_11_3 = {result[108*word_length*2-1 -: word_length*2]};
assign pixels_12_3 = {result[109*word_length*2-1 -: word_length*2]};
assign pixels_13_3 = {result[110*word_length*2-1 -: word_length*2]};
assign pixels_14_3 = {result[111*word_length*2-1 -: word_length*2]};
assign pixels_15_3 = {result[112*word_length*2-1 -: word_length*2]};
assign pixels_16_3 = {result[113*word_length*2-1 -: word_length*2]};
assign pixels_17_3 = {result[114*word_length*2-1 -: word_length*2]};
assign pixels_18_3 = {result[115*word_length*2-1 -: word_length*2]};
assign pixels_19_3 = {result[116*word_length*2-1 -: word_length*2]};
assign pixels_20_3 = {result[117*word_length*2-1 -: word_length*2]};
assign pixels_21_3 = {result[118*word_length*2-1 -: word_length*2]};
assign pixels_22_3 = {result[119*word_length*2-1 -: word_length*2]};
assign pixels_23_3 = {result[120*word_length*2-1 -: word_length*2]};
assign pixels_24_3 = {result[121*word_length*2-1 -: word_length*2]};
assign pixels_25_3 = {result[122*word_length*2-1 -: word_length*2]};
assign pixels_26_3 = {result[123*word_length*2-1 -: word_length*2]};
assign pixels_27_3 = {result[124*word_length*2-1 -: word_length*2]};
assign pixels_28_3 = {result[125*word_length*2-1 -: word_length*2]};
assign pixels_29_3 = {result[126*word_length*2-1 -: word_length*2]};
assign pixels_30_3 = {result[127*word_length*2-1 -: word_length*2]};
assign pixels_31_3 = {result[128*word_length*2-1 -: word_length*2]};
assign pixels_0_4 = {result[129*word_length*2-1 -: word_length*2]};
assign pixels_1_4 = {result[130*word_length*2-1 -: word_length*2]};
assign pixels_2_4 = {result[131*word_length*2-1 -: word_length*2]};
assign pixels_3_4 = {result[132*word_length*2-1 -: word_length*2]};
assign pixels_4_4 = {result[133*word_length*2-1 -: word_length*2]};
assign pixels_5_4 = {result[134*word_length*2-1 -: word_length*2]};
assign pixels_6_4 = {result[135*word_length*2-1 -: word_length*2]};
assign pixels_7_4 = {result[136*word_length*2-1 -: word_length*2]};
assign pixels_8_4 = {result[137*word_length*2-1 -: word_length*2]};
assign pixels_9_4 = {result[138*word_length*2-1 -: word_length*2]};
assign pixels_10_4 = {result[139*word_length*2-1 -: word_length*2]};
assign pixels_11_4 = {result[140*word_length*2-1 -: word_length*2]};
assign pixels_12_4 = {result[141*word_length*2-1 -: word_length*2]};
assign pixels_13_4 = {result[142*word_length*2-1 -: word_length*2]};
assign pixels_14_4 = {result[143*word_length*2-1 -: word_length*2]};
assign pixels_15_4 = {result[144*word_length*2-1 -: word_length*2]};
assign pixels_16_4 = {result[145*word_length*2-1 -: word_length*2]};
assign pixels_17_4 = {result[146*word_length*2-1 -: word_length*2]};
assign pixels_18_4 = {result[147*word_length*2-1 -: word_length*2]};
assign pixels_19_4 = {result[148*word_length*2-1 -: word_length*2]};
assign pixels_20_4 = {result[149*word_length*2-1 -: word_length*2]};
assign pixels_21_4 = {result[150*word_length*2-1 -: word_length*2]};
assign pixels_22_4 = {result[151*word_length*2-1 -: word_length*2]};
assign pixels_23_4 = {result[152*word_length*2-1 -: word_length*2]};
assign pixels_24_4 = {result[153*word_length*2-1 -: word_length*2]};
assign pixels_25_4 = {result[154*word_length*2-1 -: word_length*2]};
assign pixels_26_4 = {result[155*word_length*2-1 -: word_length*2]};
assign pixels_27_4 = {result[156*word_length*2-1 -: word_length*2]};
assign pixels_28_4 = {result[157*word_length*2-1 -: word_length*2]};
assign pixels_29_4 = {result[158*word_length*2-1 -: word_length*2]};
assign pixels_30_4 = {result[159*word_length*2-1 -: word_length*2]};
assign pixels_31_4 = {result[160*word_length*2-1 -: word_length*2]};
assign pixels_0_5 = {result[161*word_length*2-1 -: word_length*2]};
assign pixels_1_5 = {result[162*word_length*2-1 -: word_length*2]};
assign pixels_2_5 = {result[163*word_length*2-1 -: word_length*2]};
assign pixels_3_5 = {result[164*word_length*2-1 -: word_length*2]};
assign pixels_4_5 = {result[165*word_length*2-1 -: word_length*2]};
assign pixels_5_5 = {result[166*word_length*2-1 -: word_length*2]};
assign pixels_6_5 = {result[167*word_length*2-1 -: word_length*2]};
assign pixels_7_5 = {result[168*word_length*2-1 -: word_length*2]};
assign pixels_8_5 = {result[169*word_length*2-1 -: word_length*2]};
assign pixels_9_5 = {result[170*word_length*2-1 -: word_length*2]};
assign pixels_10_5 = {result[171*word_length*2-1 -: word_length*2]};
assign pixels_11_5 = {result[172*word_length*2-1 -: word_length*2]};
assign pixels_12_5 = {result[173*word_length*2-1 -: word_length*2]};
assign pixels_13_5 = {result[174*word_length*2-1 -: word_length*2]};
assign pixels_14_5 = {result[175*word_length*2-1 -: word_length*2]};
assign pixels_15_5 = {result[176*word_length*2-1 -: word_length*2]};
assign pixels_16_5 = {result[177*word_length*2-1 -: word_length*2]};
assign pixels_17_5 = {result[178*word_length*2-1 -: word_length*2]};
assign pixels_18_5 = {result[179*word_length*2-1 -: word_length*2]};
assign pixels_19_5 = {result[180*word_length*2-1 -: word_length*2]};
assign pixels_20_5 = {result[181*word_length*2-1 -: word_length*2]};
assign pixels_21_5 = {result[182*word_length*2-1 -: word_length*2]};
assign pixels_22_5 = {result[183*word_length*2-1 -: word_length*2]};
assign pixels_23_5 = {result[184*word_length*2-1 -: word_length*2]};
assign pixels_24_5 = {result[185*word_length*2-1 -: word_length*2]};
assign pixels_25_5 = {result[186*word_length*2-1 -: word_length*2]};
assign pixels_26_5 = {result[187*word_length*2-1 -: word_length*2]};
assign pixels_27_5 = {result[188*word_length*2-1 -: word_length*2]};
assign pixels_28_5 = {result[189*word_length*2-1 -: word_length*2]};
assign pixels_29_5 = {result[190*word_length*2-1 -: word_length*2]};
assign pixels_30_5 = {result[191*word_length*2-1 -: word_length*2]};
assign pixels_31_5 = {result[192*word_length*2-1 -: word_length*2]};
assign pixels_0_6 = {result[193*word_length*2-1 -: word_length*2]};
assign pixels_1_6 = {result[194*word_length*2-1 -: word_length*2]};
assign pixels_2_6 = {result[195*word_length*2-1 -: word_length*2]};
assign pixels_3_6 = {result[196*word_length*2-1 -: word_length*2]};
assign pixels_4_6 = {result[197*word_length*2-1 -: word_length*2]};
assign pixels_5_6 = {result[198*word_length*2-1 -: word_length*2]};
assign pixels_6_6 = {result[199*word_length*2-1 -: word_length*2]};
assign pixels_7_6 = {result[200*word_length*2-1 -: word_length*2]};
assign pixels_8_6 = {result[201*word_length*2-1 -: word_length*2]};
assign pixels_9_6 = {result[202*word_length*2-1 -: word_length*2]};
assign pixels_10_6 = {result[203*word_length*2-1 -: word_length*2]};
assign pixels_11_6 = {result[204*word_length*2-1 -: word_length*2]};
assign pixels_12_6 = {result[205*word_length*2-1 -: word_length*2]};
assign pixels_13_6 = {result[206*word_length*2-1 -: word_length*2]};
assign pixels_14_6 = {result[207*word_length*2-1 -: word_length*2]};
assign pixels_15_6 = {result[208*word_length*2-1 -: word_length*2]};
assign pixels_16_6 = {result[209*word_length*2-1 -: word_length*2]};
assign pixels_17_6 = {result[210*word_length*2-1 -: word_length*2]};
assign pixels_18_6 = {result[211*word_length*2-1 -: word_length*2]};
assign pixels_19_6 = {result[212*word_length*2-1 -: word_length*2]};
assign pixels_20_6 = {result[213*word_length*2-1 -: word_length*2]};
assign pixels_21_6 = {result[214*word_length*2-1 -: word_length*2]};
assign pixels_22_6 = {result[215*word_length*2-1 -: word_length*2]};
assign pixels_23_6 = {result[216*word_length*2-1 -: word_length*2]};
assign pixels_24_6 = {result[217*word_length*2-1 -: word_length*2]};
assign pixels_25_6 = {result[218*word_length*2-1 -: word_length*2]};
assign pixels_26_6 = {result[219*word_length*2-1 -: word_length*2]};
assign pixels_27_6 = {result[220*word_length*2-1 -: word_length*2]};
assign pixels_28_6 = {result[221*word_length*2-1 -: word_length*2]};
assign pixels_29_6 = {result[222*word_length*2-1 -: word_length*2]};
assign pixels_30_6 = {result[223*word_length*2-1 -: word_length*2]};
assign pixels_31_6 = {result[224*word_length*2-1 -: word_length*2]};
assign pixels_0_7 = {result[225*word_length*2-1 -: word_length*2]};
assign pixels_1_7 = {result[226*word_length*2-1 -: word_length*2]};
assign pixels_2_7 = {result[227*word_length*2-1 -: word_length*2]};
assign pixels_3_7 = {result[228*word_length*2-1 -: word_length*2]};
assign pixels_4_7 = {result[229*word_length*2-1 -: word_length*2]};
assign pixels_5_7 = {result[230*word_length*2-1 -: word_length*2]};
assign pixels_6_7 = {result[231*word_length*2-1 -: word_length*2]};
assign pixels_7_7 = {result[232*word_length*2-1 -: word_length*2]};
assign pixels_8_7 = {result[233*word_length*2-1 -: word_length*2]};
assign pixels_9_7 = {result[234*word_length*2-1 -: word_length*2]};
assign pixels_10_7 = {result[235*word_length*2-1 -: word_length*2]};
assign pixels_11_7 = {result[236*word_length*2-1 -: word_length*2]};
assign pixels_12_7 = {result[237*word_length*2-1 -: word_length*2]};
assign pixels_13_7 = {result[238*word_length*2-1 -: word_length*2]};
assign pixels_14_7 = {result[239*word_length*2-1 -: word_length*2]};
assign pixels_15_7 = {result[240*word_length*2-1 -: word_length*2]};
assign pixels_16_7 = {result[241*word_length*2-1 -: word_length*2]};
assign pixels_17_7 = {result[242*word_length*2-1 -: word_length*2]};
assign pixels_18_7 = {result[243*word_length*2-1 -: word_length*2]};
assign pixels_19_7 = {result[244*word_length*2-1 -: word_length*2]};
assign pixels_20_7 = {result[245*word_length*2-1 -: word_length*2]};
assign pixels_21_7 = {result[246*word_length*2-1 -: word_length*2]};
assign pixels_22_7 = {result[247*word_length*2-1 -: word_length*2]};
assign pixels_23_7 = {result[248*word_length*2-1 -: word_length*2]};
assign pixels_24_7 = {result[249*word_length*2-1 -: word_length*2]};
assign pixels_25_7 = {result[250*word_length*2-1 -: word_length*2]};
assign pixels_26_7 = {result[251*word_length*2-1 -: word_length*2]};
assign pixels_27_7 = {result[252*word_length*2-1 -: word_length*2]};
assign pixels_28_7 = {result[253*word_length*2-1 -: word_length*2]};
assign pixels_29_7 = {result[254*word_length*2-1 -: word_length*2]};
assign pixels_30_7 = {result[255*word_length*2-1 -: word_length*2]};
assign pixels_31_7 = {result[256*word_length*2-1 -: word_length*2]};
assign pixels_0_8 = {result[257*word_length*2-1 -: word_length*2]};
assign pixels_1_8 = {result[258*word_length*2-1 -: word_length*2]};
assign pixels_2_8 = {result[259*word_length*2-1 -: word_length*2]};
assign pixels_3_8 = {result[260*word_length*2-1 -: word_length*2]};
assign pixels_4_8 = {result[261*word_length*2-1 -: word_length*2]};
assign pixels_5_8 = {result[262*word_length*2-1 -: word_length*2]};
assign pixels_6_8 = {result[263*word_length*2-1 -: word_length*2]};
assign pixels_7_8 = {result[264*word_length*2-1 -: word_length*2]};
assign pixels_8_8 = {result[265*word_length*2-1 -: word_length*2]};
assign pixels_9_8 = {result[266*word_length*2-1 -: word_length*2]};
assign pixels_10_8 = {result[267*word_length*2-1 -: word_length*2]};
assign pixels_11_8 = {result[268*word_length*2-1 -: word_length*2]};
assign pixels_12_8 = {result[269*word_length*2-1 -: word_length*2]};
assign pixels_13_8 = {result[270*word_length*2-1 -: word_length*2]};
assign pixels_14_8 = {result[271*word_length*2-1 -: word_length*2]};
assign pixels_15_8 = {result[272*word_length*2-1 -: word_length*2]};
assign pixels_16_8 = {result[273*word_length*2-1 -: word_length*2]};
assign pixels_17_8 = {result[274*word_length*2-1 -: word_length*2]};
assign pixels_18_8 = {result[275*word_length*2-1 -: word_length*2]};
assign pixels_19_8 = {result[276*word_length*2-1 -: word_length*2]};
assign pixels_20_8 = {result[277*word_length*2-1 -: word_length*2]};
assign pixels_21_8 = {result[278*word_length*2-1 -: word_length*2]};
assign pixels_22_8 = {result[279*word_length*2-1 -: word_length*2]};
assign pixels_23_8 = {result[280*word_length*2-1 -: word_length*2]};
assign pixels_24_8 = {result[281*word_length*2-1 -: word_length*2]};
assign pixels_25_8 = {result[282*word_length*2-1 -: word_length*2]};
assign pixels_26_8 = {result[283*word_length*2-1 -: word_length*2]};
assign pixels_27_8 = {result[284*word_length*2-1 -: word_length*2]};
assign pixels_28_8 = {result[285*word_length*2-1 -: word_length*2]};
assign pixels_29_8 = {result[286*word_length*2-1 -: word_length*2]};
assign pixels_30_8 = {result[287*word_length*2-1 -: word_length*2]};
assign pixels_31_8 = {result[288*word_length*2-1 -: word_length*2]};
assign pixels_0_9 = {result[289*word_length*2-1 -: word_length*2]};
assign pixels_1_9 = {result[290*word_length*2-1 -: word_length*2]};
assign pixels_2_9 = {result[291*word_length*2-1 -: word_length*2]};
assign pixels_3_9 = {result[292*word_length*2-1 -: word_length*2]};
assign pixels_4_9 = {result[293*word_length*2-1 -: word_length*2]};
assign pixels_5_9 = {result[294*word_length*2-1 -: word_length*2]};
assign pixels_6_9 = {result[295*word_length*2-1 -: word_length*2]};
assign pixels_7_9 = {result[296*word_length*2-1 -: word_length*2]};
assign pixels_8_9 = {result[297*word_length*2-1 -: word_length*2]};
assign pixels_9_9 = {result[298*word_length*2-1 -: word_length*2]};
assign pixels_10_9 = {result[299*word_length*2-1 -: word_length*2]};
assign pixels_11_9 = {result[300*word_length*2-1 -: word_length*2]};
assign pixels_12_9 = {result[301*word_length*2-1 -: word_length*2]};
assign pixels_13_9 = {result[302*word_length*2-1 -: word_length*2]};
assign pixels_14_9 = {result[303*word_length*2-1 -: word_length*2]};
assign pixels_15_9 = {result[304*word_length*2-1 -: word_length*2]};
assign pixels_16_9 = {result[305*word_length*2-1 -: word_length*2]};
assign pixels_17_9 = {result[306*word_length*2-1 -: word_length*2]};
assign pixels_18_9 = {result[307*word_length*2-1 -: word_length*2]};
assign pixels_19_9 = {result[308*word_length*2-1 -: word_length*2]};
assign pixels_20_9 = {result[309*word_length*2-1 -: word_length*2]};
assign pixels_21_9 = {result[310*word_length*2-1 -: word_length*2]};
assign pixels_22_9 = {result[311*word_length*2-1 -: word_length*2]};
assign pixels_23_9 = {result[312*word_length*2-1 -: word_length*2]};
assign pixels_24_9 = {result[313*word_length*2-1 -: word_length*2]};
assign pixels_25_9 = {result[314*word_length*2-1 -: word_length*2]};
assign pixels_26_9 = {result[315*word_length*2-1 -: word_length*2]};
assign pixels_27_9 = {result[316*word_length*2-1 -: word_length*2]};
assign pixels_28_9 = {result[317*word_length*2-1 -: word_length*2]};
assign pixels_29_9 = {result[318*word_length*2-1 -: word_length*2]};
assign pixels_30_9 = {result[319*word_length*2-1 -: word_length*2]};
assign pixels_31_9 = {result[320*word_length*2-1 -: word_length*2]};
assign pixels_0_10 = {result[321*word_length*2-1 -: word_length*2]};
assign pixels_1_10 = {result[322*word_length*2-1 -: word_length*2]};
assign pixels_2_10 = {result[323*word_length*2-1 -: word_length*2]};
assign pixels_3_10 = {result[324*word_length*2-1 -: word_length*2]};
assign pixels_4_10 = {result[325*word_length*2-1 -: word_length*2]};
assign pixels_5_10 = {result[326*word_length*2-1 -: word_length*2]};
assign pixels_6_10 = {result[327*word_length*2-1 -: word_length*2]};
assign pixels_7_10 = {result[328*word_length*2-1 -: word_length*2]};
assign pixels_8_10 = {result[329*word_length*2-1 -: word_length*2]};
assign pixels_9_10 = {result[330*word_length*2-1 -: word_length*2]};
assign pixels_10_10 = {result[331*word_length*2-1 -: word_length*2]};
assign pixels_11_10 = {result[332*word_length*2-1 -: word_length*2]};
assign pixels_12_10 = {result[333*word_length*2-1 -: word_length*2]};
assign pixels_13_10 = {result[334*word_length*2-1 -: word_length*2]};
assign pixels_14_10 = {result[335*word_length*2-1 -: word_length*2]};
assign pixels_15_10 = {result[336*word_length*2-1 -: word_length*2]};
assign pixels_16_10 = {result[337*word_length*2-1 -: word_length*2]};
assign pixels_17_10 = {result[338*word_length*2-1 -: word_length*2]};
assign pixels_18_10 = {result[339*word_length*2-1 -: word_length*2]};
assign pixels_19_10 = {result[340*word_length*2-1 -: word_length*2]};
assign pixels_20_10 = {result[341*word_length*2-1 -: word_length*2]};
assign pixels_21_10 = {result[342*word_length*2-1 -: word_length*2]};
assign pixels_22_10 = {result[343*word_length*2-1 -: word_length*2]};
assign pixels_23_10 = {result[344*word_length*2-1 -: word_length*2]};
assign pixels_24_10 = {result[345*word_length*2-1 -: word_length*2]};
assign pixels_25_10 = {result[346*word_length*2-1 -: word_length*2]};
assign pixels_26_10 = {result[347*word_length*2-1 -: word_length*2]};
assign pixels_27_10 = {result[348*word_length*2-1 -: word_length*2]};
assign pixels_28_10 = {result[349*word_length*2-1 -: word_length*2]};
assign pixels_29_10 = {result[350*word_length*2-1 -: word_length*2]};
assign pixels_30_10 = {result[351*word_length*2-1 -: word_length*2]};
assign pixels_31_10 = {result[352*word_length*2-1 -: word_length*2]};
assign pixels_0_11 = {result[353*word_length*2-1 -: word_length*2]};
assign pixels_1_11 = {result[354*word_length*2-1 -: word_length*2]};
assign pixels_2_11 = {result[355*word_length*2-1 -: word_length*2]};
assign pixels_3_11 = {result[356*word_length*2-1 -: word_length*2]};
assign pixels_4_11 = {result[357*word_length*2-1 -: word_length*2]};
assign pixels_5_11 = {result[358*word_length*2-1 -: word_length*2]};
assign pixels_6_11 = {result[359*word_length*2-1 -: word_length*2]};
assign pixels_7_11 = {result[360*word_length*2-1 -: word_length*2]};
assign pixels_8_11 = {result[361*word_length*2-1 -: word_length*2]};
assign pixels_9_11 = {result[362*word_length*2-1 -: word_length*2]};
assign pixels_10_11 = {result[363*word_length*2-1 -: word_length*2]};
assign pixels_11_11 = {result[364*word_length*2-1 -: word_length*2]};
assign pixels_12_11 = {result[365*word_length*2-1 -: word_length*2]};
assign pixels_13_11 = {result[366*word_length*2-1 -: word_length*2]};
assign pixels_14_11 = {result[367*word_length*2-1 -: word_length*2]};
assign pixels_15_11 = {result[368*word_length*2-1 -: word_length*2]};
assign pixels_16_11 = {result[369*word_length*2-1 -: word_length*2]};
assign pixels_17_11 = {result[370*word_length*2-1 -: word_length*2]};
assign pixels_18_11 = {result[371*word_length*2-1 -: word_length*2]};
assign pixels_19_11 = {result[372*word_length*2-1 -: word_length*2]};
assign pixels_20_11 = {result[373*word_length*2-1 -: word_length*2]};
assign pixels_21_11 = {result[374*word_length*2-1 -: word_length*2]};
assign pixels_22_11 = {result[375*word_length*2-1 -: word_length*2]};
assign pixels_23_11 = {result[376*word_length*2-1 -: word_length*2]};
assign pixels_24_11 = {result[377*word_length*2-1 -: word_length*2]};
assign pixels_25_11 = {result[378*word_length*2-1 -: word_length*2]};
assign pixels_26_11 = {result[379*word_length*2-1 -: word_length*2]};
assign pixels_27_11 = {result[380*word_length*2-1 -: word_length*2]};
assign pixels_28_11 = {result[381*word_length*2-1 -: word_length*2]};
assign pixels_29_11 = {result[382*word_length*2-1 -: word_length*2]};
assign pixels_30_11 = {result[383*word_length*2-1 -: word_length*2]};
assign pixels_31_11 = {result[384*word_length*2-1 -: word_length*2]};
assign pixels_0_12 = {result[385*word_length*2-1 -: word_length*2]};
assign pixels_1_12 = {result[386*word_length*2-1 -: word_length*2]};
assign pixels_2_12 = {result[387*word_length*2-1 -: word_length*2]};
assign pixels_3_12 = {result[388*word_length*2-1 -: word_length*2]};
assign pixels_4_12 = {result[389*word_length*2-1 -: word_length*2]};
assign pixels_5_12 = {result[390*word_length*2-1 -: word_length*2]};
assign pixels_6_12 = {result[391*word_length*2-1 -: word_length*2]};
assign pixels_7_12 = {result[392*word_length*2-1 -: word_length*2]};
assign pixels_8_12 = {result[393*word_length*2-1 -: word_length*2]};
assign pixels_9_12 = {result[394*word_length*2-1 -: word_length*2]};
assign pixels_10_12 = {result[395*word_length*2-1 -: word_length*2]};
assign pixels_11_12 = {result[396*word_length*2-1 -: word_length*2]};
assign pixels_12_12 = {result[397*word_length*2-1 -: word_length*2]};
assign pixels_13_12 = {result[398*word_length*2-1 -: word_length*2]};
assign pixels_14_12 = {result[399*word_length*2-1 -: word_length*2]};
assign pixels_15_12 = {result[400*word_length*2-1 -: word_length*2]};
assign pixels_16_12 = {result[401*word_length*2-1 -: word_length*2]};
assign pixels_17_12 = {result[402*word_length*2-1 -: word_length*2]};
assign pixels_18_12 = {result[403*word_length*2-1 -: word_length*2]};
assign pixels_19_12 = {result[404*word_length*2-1 -: word_length*2]};
assign pixels_20_12 = {result[405*word_length*2-1 -: word_length*2]};
assign pixels_21_12 = {result[406*word_length*2-1 -: word_length*2]};
assign pixels_22_12 = {result[407*word_length*2-1 -: word_length*2]};
assign pixels_23_12 = {result[408*word_length*2-1 -: word_length*2]};
assign pixels_24_12 = {result[409*word_length*2-1 -: word_length*2]};
assign pixels_25_12 = {result[410*word_length*2-1 -: word_length*2]};
assign pixels_26_12 = {result[411*word_length*2-1 -: word_length*2]};
assign pixels_27_12 = {result[412*word_length*2-1 -: word_length*2]};
assign pixels_28_12 = {result[413*word_length*2-1 -: word_length*2]};
assign pixels_29_12 = {result[414*word_length*2-1 -: word_length*2]};
assign pixels_30_12 = {result[415*word_length*2-1 -: word_length*2]};
assign pixels_31_12 = {result[416*word_length*2-1 -: word_length*2]};
assign pixels_0_13 = {result[417*word_length*2-1 -: word_length*2]};
assign pixels_1_13 = {result[418*word_length*2-1 -: word_length*2]};
assign pixels_2_13 = {result[419*word_length*2-1 -: word_length*2]};
assign pixels_3_13 = {result[420*word_length*2-1 -: word_length*2]};
assign pixels_4_13 = {result[421*word_length*2-1 -: word_length*2]};
assign pixels_5_13 = {result[422*word_length*2-1 -: word_length*2]};
assign pixels_6_13 = {result[423*word_length*2-1 -: word_length*2]};
assign pixels_7_13 = {result[424*word_length*2-1 -: word_length*2]};
assign pixels_8_13 = {result[425*word_length*2-1 -: word_length*2]};
assign pixels_9_13 = {result[426*word_length*2-1 -: word_length*2]};
assign pixels_10_13 = {result[427*word_length*2-1 -: word_length*2]};
assign pixels_11_13 = {result[428*word_length*2-1 -: word_length*2]};
assign pixels_12_13 = {result[429*word_length*2-1 -: word_length*2]};
assign pixels_13_13 = {result[430*word_length*2-1 -: word_length*2]};
assign pixels_14_13 = {result[431*word_length*2-1 -: word_length*2]};
assign pixels_15_13 = {result[432*word_length*2-1 -: word_length*2]};
assign pixels_16_13 = {result[433*word_length*2-1 -: word_length*2]};
assign pixels_17_13 = {result[434*word_length*2-1 -: word_length*2]};
assign pixels_18_13 = {result[435*word_length*2-1 -: word_length*2]};
assign pixels_19_13 = {result[436*word_length*2-1 -: word_length*2]};
assign pixels_20_13 = {result[437*word_length*2-1 -: word_length*2]};
assign pixels_21_13 = {result[438*word_length*2-1 -: word_length*2]};
assign pixels_22_13 = {result[439*word_length*2-1 -: word_length*2]};
assign pixels_23_13 = {result[440*word_length*2-1 -: word_length*2]};
assign pixels_24_13 = {result[441*word_length*2-1 -: word_length*2]};
assign pixels_25_13 = {result[442*word_length*2-1 -: word_length*2]};
assign pixels_26_13 = {result[443*word_length*2-1 -: word_length*2]};
assign pixels_27_13 = {result[444*word_length*2-1 -: word_length*2]};
assign pixels_28_13 = {result[445*word_length*2-1 -: word_length*2]};
assign pixels_29_13 = {result[446*word_length*2-1 -: word_length*2]};
assign pixels_30_13 = {result[447*word_length*2-1 -: word_length*2]};
assign pixels_31_13 = {result[448*word_length*2-1 -: word_length*2]};
assign pixels_0_14 = {result[449*word_length*2-1 -: word_length*2]};
assign pixels_1_14 = {result[450*word_length*2-1 -: word_length*2]};
assign pixels_2_14 = {result[451*word_length*2-1 -: word_length*2]};
assign pixels_3_14 = {result[452*word_length*2-1 -: word_length*2]};
assign pixels_4_14 = {result[453*word_length*2-1 -: word_length*2]};
assign pixels_5_14 = {result[454*word_length*2-1 -: word_length*2]};
assign pixels_6_14 = {result[455*word_length*2-1 -: word_length*2]};
assign pixels_7_14 = {result[456*word_length*2-1 -: word_length*2]};
assign pixels_8_14 = {result[457*word_length*2-1 -: word_length*2]};
assign pixels_9_14 = {result[458*word_length*2-1 -: word_length*2]};
assign pixels_10_14 = {result[459*word_length*2-1 -: word_length*2]};
assign pixels_11_14 = {result[460*word_length*2-1 -: word_length*2]};
assign pixels_12_14 = {result[461*word_length*2-1 -: word_length*2]};
assign pixels_13_14 = {result[462*word_length*2-1 -: word_length*2]};
assign pixels_14_14 = {result[463*word_length*2-1 -: word_length*2]};
assign pixels_15_14 = {result[464*word_length*2-1 -: word_length*2]};
assign pixels_16_14 = {result[465*word_length*2-1 -: word_length*2]};
assign pixels_17_14 = {result[466*word_length*2-1 -: word_length*2]};
assign pixels_18_14 = {result[467*word_length*2-1 -: word_length*2]};
assign pixels_19_14 = {result[468*word_length*2-1 -: word_length*2]};
assign pixels_20_14 = {result[469*word_length*2-1 -: word_length*2]};
assign pixels_21_14 = {result[470*word_length*2-1 -: word_length*2]};
assign pixels_22_14 = {result[471*word_length*2-1 -: word_length*2]};
assign pixels_23_14 = {result[472*word_length*2-1 -: word_length*2]};
assign pixels_24_14 = {result[473*word_length*2-1 -: word_length*2]};
assign pixels_25_14 = {result[474*word_length*2-1 -: word_length*2]};
assign pixels_26_14 = {result[475*word_length*2-1 -: word_length*2]};
assign pixels_27_14 = {result[476*word_length*2-1 -: word_length*2]};
assign pixels_28_14 = {result[477*word_length*2-1 -: word_length*2]};
assign pixels_29_14 = {result[478*word_length*2-1 -: word_length*2]};
assign pixels_30_14 = {result[479*word_length*2-1 -: word_length*2]};
assign pixels_31_14 = {result[480*word_length*2-1 -: word_length*2]};
assign pixels_0_15 = {result[481*word_length*2-1 -: word_length*2]};
assign pixels_1_15 = {result[482*word_length*2-1 -: word_length*2]};
assign pixels_2_15 = {result[483*word_length*2-1 -: word_length*2]};
assign pixels_3_15 = {result[484*word_length*2-1 -: word_length*2]};
assign pixels_4_15 = {result[485*word_length*2-1 -: word_length*2]};
assign pixels_5_15 = {result[486*word_length*2-1 -: word_length*2]};
assign pixels_6_15 = {result[487*word_length*2-1 -: word_length*2]};
assign pixels_7_15 = {result[488*word_length*2-1 -: word_length*2]};
assign pixels_8_15 = {result[489*word_length*2-1 -: word_length*2]};
assign pixels_9_15 = {result[490*word_length*2-1 -: word_length*2]};
assign pixels_10_15 = {result[491*word_length*2-1 -: word_length*2]};
assign pixels_11_15 = {result[492*word_length*2-1 -: word_length*2]};
assign pixels_12_15 = {result[493*word_length*2-1 -: word_length*2]};
assign pixels_13_15 = {result[494*word_length*2-1 -: word_length*2]};
assign pixels_14_15 = {result[495*word_length*2-1 -: word_length*2]};
assign pixels_15_15 = {result[496*word_length*2-1 -: word_length*2]};
assign pixels_16_15 = {result[497*word_length*2-1 -: word_length*2]};
assign pixels_17_15 = {result[498*word_length*2-1 -: word_length*2]};
assign pixels_18_15 = {result[499*word_length*2-1 -: word_length*2]};
assign pixels_19_15 = {result[500*word_length*2-1 -: word_length*2]};
assign pixels_20_15 = {result[501*word_length*2-1 -: word_length*2]};
assign pixels_21_15 = {result[502*word_length*2-1 -: word_length*2]};
assign pixels_22_15 = {result[503*word_length*2-1 -: word_length*2]};
assign pixels_23_15 = {result[504*word_length*2-1 -: word_length*2]};
assign pixels_24_15 = {result[505*word_length*2-1 -: word_length*2]};
assign pixels_25_15 = {result[506*word_length*2-1 -: word_length*2]};
assign pixels_26_15 = {result[507*word_length*2-1 -: word_length*2]};
assign pixels_27_15 = {result[508*word_length*2-1 -: word_length*2]};
assign pixels_28_15 = {result[509*word_length*2-1 -: word_length*2]};
assign pixels_29_15 = {result[510*word_length*2-1 -: word_length*2]};
assign pixels_30_15 = {result[511*word_length*2-1 -: word_length*2]};
assign pixels_31_15 = {result[512*word_length*2-1 -: word_length*2]};
assign pixels_0_16 = {result[513*word_length*2-1 -: word_length*2]};
assign pixels_1_16 = {result[514*word_length*2-1 -: word_length*2]};
assign pixels_2_16 = {result[515*word_length*2-1 -: word_length*2]};
assign pixels_3_16 = {result[516*word_length*2-1 -: word_length*2]};
assign pixels_4_16 = {result[517*word_length*2-1 -: word_length*2]};
assign pixels_5_16 = {result[518*word_length*2-1 -: word_length*2]};
assign pixels_6_16 = {result[519*word_length*2-1 -: word_length*2]};
assign pixels_7_16 = {result[520*word_length*2-1 -: word_length*2]};
assign pixels_8_16 = {result[521*word_length*2-1 -: word_length*2]};
assign pixels_9_16 = {result[522*word_length*2-1 -: word_length*2]};
assign pixels_10_16 = {result[523*word_length*2-1 -: word_length*2]};
assign pixels_11_16 = {result[524*word_length*2-1 -: word_length*2]};
assign pixels_12_16 = {result[525*word_length*2-1 -: word_length*2]};
assign pixels_13_16 = {result[526*word_length*2-1 -: word_length*2]};
assign pixels_14_16 = {result[527*word_length*2-1 -: word_length*2]};
assign pixels_15_16 = {result[528*word_length*2-1 -: word_length*2]};
assign pixels_16_16 = {result[529*word_length*2-1 -: word_length*2]};
assign pixels_17_16 = {result[530*word_length*2-1 -: word_length*2]};
assign pixels_18_16 = {result[531*word_length*2-1 -: word_length*2]};
assign pixels_19_16 = {result[532*word_length*2-1 -: word_length*2]};
assign pixels_20_16 = {result[533*word_length*2-1 -: word_length*2]};
assign pixels_21_16 = {result[534*word_length*2-1 -: word_length*2]};
assign pixels_22_16 = {result[535*word_length*2-1 -: word_length*2]};
assign pixels_23_16 = {result[536*word_length*2-1 -: word_length*2]};
assign pixels_24_16 = {result[537*word_length*2-1 -: word_length*2]};
assign pixels_25_16 = {result[538*word_length*2-1 -: word_length*2]};
assign pixels_26_16 = {result[539*word_length*2-1 -: word_length*2]};
assign pixels_27_16 = {result[540*word_length*2-1 -: word_length*2]};
assign pixels_28_16 = {result[541*word_length*2-1 -: word_length*2]};
assign pixels_29_16 = {result[542*word_length*2-1 -: word_length*2]};
assign pixels_30_16 = {result[543*word_length*2-1 -: word_length*2]};
assign pixels_31_16 = {result[544*word_length*2-1 -: word_length*2]};
assign pixels_0_17 = {result[545*word_length*2-1 -: word_length*2]};
assign pixels_1_17 = {result[546*word_length*2-1 -: word_length*2]};
assign pixels_2_17 = {result[547*word_length*2-1 -: word_length*2]};
assign pixels_3_17 = {result[548*word_length*2-1 -: word_length*2]};
assign pixels_4_17 = {result[549*word_length*2-1 -: word_length*2]};
assign pixels_5_17 = {result[550*word_length*2-1 -: word_length*2]};
assign pixels_6_17 = {result[551*word_length*2-1 -: word_length*2]};
assign pixels_7_17 = {result[552*word_length*2-1 -: word_length*2]};
assign pixels_8_17 = {result[553*word_length*2-1 -: word_length*2]};
assign pixels_9_17 = {result[554*word_length*2-1 -: word_length*2]};
assign pixels_10_17 = {result[555*word_length*2-1 -: word_length*2]};
assign pixels_11_17 = {result[556*word_length*2-1 -: word_length*2]};
assign pixels_12_17 = {result[557*word_length*2-1 -: word_length*2]};
assign pixels_13_17 = {result[558*word_length*2-1 -: word_length*2]};
assign pixels_14_17 = {result[559*word_length*2-1 -: word_length*2]};
assign pixels_15_17 = {result[560*word_length*2-1 -: word_length*2]};
assign pixels_16_17 = {result[561*word_length*2-1 -: word_length*2]};
assign pixels_17_17 = {result[562*word_length*2-1 -: word_length*2]};
assign pixels_18_17 = {result[563*word_length*2-1 -: word_length*2]};
assign pixels_19_17 = {result[564*word_length*2-1 -: word_length*2]};
assign pixels_20_17 = {result[565*word_length*2-1 -: word_length*2]};
assign pixels_21_17 = {result[566*word_length*2-1 -: word_length*2]};
assign pixels_22_17 = {result[567*word_length*2-1 -: word_length*2]};
assign pixels_23_17 = {result[568*word_length*2-1 -: word_length*2]};
assign pixels_24_17 = {result[569*word_length*2-1 -: word_length*2]};
assign pixels_25_17 = {result[570*word_length*2-1 -: word_length*2]};
assign pixels_26_17 = {result[571*word_length*2-1 -: word_length*2]};
assign pixels_27_17 = {result[572*word_length*2-1 -: word_length*2]};
assign pixels_28_17 = {result[573*word_length*2-1 -: word_length*2]};
assign pixels_29_17 = {result[574*word_length*2-1 -: word_length*2]};
assign pixels_30_17 = {result[575*word_length*2-1 -: word_length*2]};
assign pixels_31_17 = {result[576*word_length*2-1 -: word_length*2]};
assign pixels_0_18 = {result[577*word_length*2-1 -: word_length*2]};
assign pixels_1_18 = {result[578*word_length*2-1 -: word_length*2]};
assign pixels_2_18 = {result[579*word_length*2-1 -: word_length*2]};
assign pixels_3_18 = {result[580*word_length*2-1 -: word_length*2]};
assign pixels_4_18 = {result[581*word_length*2-1 -: word_length*2]};
assign pixels_5_18 = {result[582*word_length*2-1 -: word_length*2]};
assign pixels_6_18 = {result[583*word_length*2-1 -: word_length*2]};
assign pixels_7_18 = {result[584*word_length*2-1 -: word_length*2]};
assign pixels_8_18 = {result[585*word_length*2-1 -: word_length*2]};
assign pixels_9_18 = {result[586*word_length*2-1 -: word_length*2]};
assign pixels_10_18 = {result[587*word_length*2-1 -: word_length*2]};
assign pixels_11_18 = {result[588*word_length*2-1 -: word_length*2]};
assign pixels_12_18 = {result[589*word_length*2-1 -: word_length*2]};
assign pixels_13_18 = {result[590*word_length*2-1 -: word_length*2]};
assign pixels_14_18 = {result[591*word_length*2-1 -: word_length*2]};
assign pixels_15_18 = {result[592*word_length*2-1 -: word_length*2]};
assign pixels_16_18 = {result[593*word_length*2-1 -: word_length*2]};
assign pixels_17_18 = {result[594*word_length*2-1 -: word_length*2]};
assign pixels_18_18 = {result[595*word_length*2-1 -: word_length*2]};
assign pixels_19_18 = {result[596*word_length*2-1 -: word_length*2]};
assign pixels_20_18 = {result[597*word_length*2-1 -: word_length*2]};
assign pixels_21_18 = {result[598*word_length*2-1 -: word_length*2]};
assign pixels_22_18 = {result[599*word_length*2-1 -: word_length*2]};
assign pixels_23_18 = {result[600*word_length*2-1 -: word_length*2]};
assign pixels_24_18 = {result[601*word_length*2-1 -: word_length*2]};
assign pixels_25_18 = {result[602*word_length*2-1 -: word_length*2]};
assign pixels_26_18 = {result[603*word_length*2-1 -: word_length*2]};
assign pixels_27_18 = {result[604*word_length*2-1 -: word_length*2]};
assign pixels_28_18 = {result[605*word_length*2-1 -: word_length*2]};
assign pixels_29_18 = {result[606*word_length*2-1 -: word_length*2]};
assign pixels_30_18 = {result[607*word_length*2-1 -: word_length*2]};
assign pixels_31_18 = {result[608*word_length*2-1 -: word_length*2]};
assign pixels_0_19 = {result[609*word_length*2-1 -: word_length*2]};
assign pixels_1_19 = {result[610*word_length*2-1 -: word_length*2]};
assign pixels_2_19 = {result[611*word_length*2-1 -: word_length*2]};
assign pixels_3_19 = {result[612*word_length*2-1 -: word_length*2]};
assign pixels_4_19 = {result[613*word_length*2-1 -: word_length*2]};
assign pixels_5_19 = {result[614*word_length*2-1 -: word_length*2]};
assign pixels_6_19 = {result[615*word_length*2-1 -: word_length*2]};
assign pixels_7_19 = {result[616*word_length*2-1 -: word_length*2]};
assign pixels_8_19 = {result[617*word_length*2-1 -: word_length*2]};
assign pixels_9_19 = {result[618*word_length*2-1 -: word_length*2]};
assign pixels_10_19 = {result[619*word_length*2-1 -: word_length*2]};
assign pixels_11_19 = {result[620*word_length*2-1 -: word_length*2]};
assign pixels_12_19 = {result[621*word_length*2-1 -: word_length*2]};
assign pixels_13_19 = {result[622*word_length*2-1 -: word_length*2]};
assign pixels_14_19 = {result[623*word_length*2-1 -: word_length*2]};
assign pixels_15_19 = {result[624*word_length*2-1 -: word_length*2]};
assign pixels_16_19 = {result[625*word_length*2-1 -: word_length*2]};
assign pixels_17_19 = {result[626*word_length*2-1 -: word_length*2]};
assign pixels_18_19 = {result[627*word_length*2-1 -: word_length*2]};
assign pixels_19_19 = {result[628*word_length*2-1 -: word_length*2]};
assign pixels_20_19 = {result[629*word_length*2-1 -: word_length*2]};
assign pixels_21_19 = {result[630*word_length*2-1 -: word_length*2]};
assign pixels_22_19 = {result[631*word_length*2-1 -: word_length*2]};
assign pixels_23_19 = {result[632*word_length*2-1 -: word_length*2]};
assign pixels_24_19 = {result[633*word_length*2-1 -: word_length*2]};
assign pixels_25_19 = {result[634*word_length*2-1 -: word_length*2]};
assign pixels_26_19 = {result[635*word_length*2-1 -: word_length*2]};
assign pixels_27_19 = {result[636*word_length*2-1 -: word_length*2]};
assign pixels_28_19 = {result[637*word_length*2-1 -: word_length*2]};
assign pixels_29_19 = {result[638*word_length*2-1 -: word_length*2]};
assign pixels_30_19 = {result[639*word_length*2-1 -: word_length*2]};
assign pixels_31_19 = {result[640*word_length*2-1 -: word_length*2]};
assign pixels_0_20 = {result[641*word_length*2-1 -: word_length*2]};
assign pixels_1_20 = {result[642*word_length*2-1 -: word_length*2]};
assign pixels_2_20 = {result[643*word_length*2-1 -: word_length*2]};
assign pixels_3_20 = {result[644*word_length*2-1 -: word_length*2]};
assign pixels_4_20 = {result[645*word_length*2-1 -: word_length*2]};
assign pixels_5_20 = {result[646*word_length*2-1 -: word_length*2]};
assign pixels_6_20 = {result[647*word_length*2-1 -: word_length*2]};
assign pixels_7_20 = {result[648*word_length*2-1 -: word_length*2]};
assign pixels_8_20 = {result[649*word_length*2-1 -: word_length*2]};
assign pixels_9_20 = {result[650*word_length*2-1 -: word_length*2]};
assign pixels_10_20 = {result[651*word_length*2-1 -: word_length*2]};
assign pixels_11_20 = {result[652*word_length*2-1 -: word_length*2]};
assign pixels_12_20 = {result[653*word_length*2-1 -: word_length*2]};
assign pixels_13_20 = {result[654*word_length*2-1 -: word_length*2]};
assign pixels_14_20 = {result[655*word_length*2-1 -: word_length*2]};
assign pixels_15_20 = {result[656*word_length*2-1 -: word_length*2]};
assign pixels_16_20 = {result[657*word_length*2-1 -: word_length*2]};
assign pixels_17_20 = {result[658*word_length*2-1 -: word_length*2]};
assign pixels_18_20 = {result[659*word_length*2-1 -: word_length*2]};
assign pixels_19_20 = {result[660*word_length*2-1 -: word_length*2]};
assign pixels_20_20 = {result[661*word_length*2-1 -: word_length*2]};
assign pixels_21_20 = {result[662*word_length*2-1 -: word_length*2]};
assign pixels_22_20 = {result[663*word_length*2-1 -: word_length*2]};
assign pixels_23_20 = {result[664*word_length*2-1 -: word_length*2]};
assign pixels_24_20 = {result[665*word_length*2-1 -: word_length*2]};
assign pixels_25_20 = {result[666*word_length*2-1 -: word_length*2]};
assign pixels_26_20 = {result[667*word_length*2-1 -: word_length*2]};
assign pixels_27_20 = {result[668*word_length*2-1 -: word_length*2]};
assign pixels_28_20 = {result[669*word_length*2-1 -: word_length*2]};
assign pixels_29_20 = {result[670*word_length*2-1 -: word_length*2]};
assign pixels_30_20 = {result[671*word_length*2-1 -: word_length*2]};
assign pixels_31_20 = {result[672*word_length*2-1 -: word_length*2]};
assign pixels_0_21 = {result[673*word_length*2-1 -: word_length*2]};
assign pixels_1_21 = {result[674*word_length*2-1 -: word_length*2]};
assign pixels_2_21 = {result[675*word_length*2-1 -: word_length*2]};
assign pixels_3_21 = {result[676*word_length*2-1 -: word_length*2]};
assign pixels_4_21 = {result[677*word_length*2-1 -: word_length*2]};
assign pixels_5_21 = {result[678*word_length*2-1 -: word_length*2]};
assign pixels_6_21 = {result[679*word_length*2-1 -: word_length*2]};
assign pixels_7_21 = {result[680*word_length*2-1 -: word_length*2]};
assign pixels_8_21 = {result[681*word_length*2-1 -: word_length*2]};
assign pixels_9_21 = {result[682*word_length*2-1 -: word_length*2]};
assign pixels_10_21 = {result[683*word_length*2-1 -: word_length*2]};
assign pixels_11_21 = {result[684*word_length*2-1 -: word_length*2]};
assign pixels_12_21 = {result[685*word_length*2-1 -: word_length*2]};
assign pixels_13_21 = {result[686*word_length*2-1 -: word_length*2]};
assign pixels_14_21 = {result[687*word_length*2-1 -: word_length*2]};
assign pixels_15_21 = {result[688*word_length*2-1 -: word_length*2]};
assign pixels_16_21 = {result[689*word_length*2-1 -: word_length*2]};
assign pixels_17_21 = {result[690*word_length*2-1 -: word_length*2]};
assign pixels_18_21 = {result[691*word_length*2-1 -: word_length*2]};
assign pixels_19_21 = {result[692*word_length*2-1 -: word_length*2]};
assign pixels_20_21 = {result[693*word_length*2-1 -: word_length*2]};
assign pixels_21_21 = {result[694*word_length*2-1 -: word_length*2]};
assign pixels_22_21 = {result[695*word_length*2-1 -: word_length*2]};
assign pixels_23_21 = {result[696*word_length*2-1 -: word_length*2]};
assign pixels_24_21 = {result[697*word_length*2-1 -: word_length*2]};
assign pixels_25_21 = {result[698*word_length*2-1 -: word_length*2]};
assign pixels_26_21 = {result[699*word_length*2-1 -: word_length*2]};
assign pixels_27_21 = {result[700*word_length*2-1 -: word_length*2]};
assign pixels_28_21 = {result[701*word_length*2-1 -: word_length*2]};
assign pixels_29_21 = {result[702*word_length*2-1 -: word_length*2]};
assign pixels_30_21 = {result[703*word_length*2-1 -: word_length*2]};
assign pixels_31_21 = {result[704*word_length*2-1 -: word_length*2]};
assign pixels_0_22 = {result[705*word_length*2-1 -: word_length*2]};
assign pixels_1_22 = {result[706*word_length*2-1 -: word_length*2]};
assign pixels_2_22 = {result[707*word_length*2-1 -: word_length*2]};
assign pixels_3_22 = {result[708*word_length*2-1 -: word_length*2]};
assign pixels_4_22 = {result[709*word_length*2-1 -: word_length*2]};
assign pixels_5_22 = {result[710*word_length*2-1 -: word_length*2]};
assign pixels_6_22 = {result[711*word_length*2-1 -: word_length*2]};
assign pixels_7_22 = {result[712*word_length*2-1 -: word_length*2]};
assign pixels_8_22 = {result[713*word_length*2-1 -: word_length*2]};
assign pixels_9_22 = {result[714*word_length*2-1 -: word_length*2]};
assign pixels_10_22 = {result[715*word_length*2-1 -: word_length*2]};
assign pixels_11_22 = {result[716*word_length*2-1 -: word_length*2]};
assign pixels_12_22 = {result[717*word_length*2-1 -: word_length*2]};
assign pixels_13_22 = {result[718*word_length*2-1 -: word_length*2]};
assign pixels_14_22 = {result[719*word_length*2-1 -: word_length*2]};
assign pixels_15_22 = {result[720*word_length*2-1 -: word_length*2]};
assign pixels_16_22 = {result[721*word_length*2-1 -: word_length*2]};
assign pixels_17_22 = {result[722*word_length*2-1 -: word_length*2]};
assign pixels_18_22 = {result[723*word_length*2-1 -: word_length*2]};
assign pixels_19_22 = {result[724*word_length*2-1 -: word_length*2]};
assign pixels_20_22 = {result[725*word_length*2-1 -: word_length*2]};
assign pixels_21_22 = {result[726*word_length*2-1 -: word_length*2]};
assign pixels_22_22 = {result[727*word_length*2-1 -: word_length*2]};
assign pixels_23_22 = {result[728*word_length*2-1 -: word_length*2]};
assign pixels_24_22 = {result[729*word_length*2-1 -: word_length*2]};
assign pixels_25_22 = {result[730*word_length*2-1 -: word_length*2]};
assign pixels_26_22 = {result[731*word_length*2-1 -: word_length*2]};
assign pixels_27_22 = {result[732*word_length*2-1 -: word_length*2]};
assign pixels_28_22 = {result[733*word_length*2-1 -: word_length*2]};
assign pixels_29_22 = {result[734*word_length*2-1 -: word_length*2]};
assign pixels_30_22 = {result[735*word_length*2-1 -: word_length*2]};
assign pixels_31_22 = {result[736*word_length*2-1 -: word_length*2]};
assign pixels_0_23 = {result[737*word_length*2-1 -: word_length*2]};
assign pixels_1_23 = {result[738*word_length*2-1 -: word_length*2]};
assign pixels_2_23 = {result[739*word_length*2-1 -: word_length*2]};
assign pixels_3_23 = {result[740*word_length*2-1 -: word_length*2]};
assign pixels_4_23 = {result[741*word_length*2-1 -: word_length*2]};
assign pixels_5_23 = {result[742*word_length*2-1 -: word_length*2]};
assign pixels_6_23 = {result[743*word_length*2-1 -: word_length*2]};
assign pixels_7_23 = {result[744*word_length*2-1 -: word_length*2]};
assign pixels_8_23 = {result[745*word_length*2-1 -: word_length*2]};
assign pixels_9_23 = {result[746*word_length*2-1 -: word_length*2]};
assign pixels_10_23 = {result[747*word_length*2-1 -: word_length*2]};
assign pixels_11_23 = {result[748*word_length*2-1 -: word_length*2]};
assign pixels_12_23 = {result[749*word_length*2-1 -: word_length*2]};
assign pixels_13_23 = {result[750*word_length*2-1 -: word_length*2]};
assign pixels_14_23 = {result[751*word_length*2-1 -: word_length*2]};
assign pixels_15_23 = {result[752*word_length*2-1 -: word_length*2]};
assign pixels_16_23 = {result[753*word_length*2-1 -: word_length*2]};
assign pixels_17_23 = {result[754*word_length*2-1 -: word_length*2]};
assign pixels_18_23 = {result[755*word_length*2-1 -: word_length*2]};
assign pixels_19_23 = {result[756*word_length*2-1 -: word_length*2]};
assign pixels_20_23 = {result[757*word_length*2-1 -: word_length*2]};
assign pixels_21_23 = {result[758*word_length*2-1 -: word_length*2]};
assign pixels_22_23 = {result[759*word_length*2-1 -: word_length*2]};
assign pixels_23_23 = {result[760*word_length*2-1 -: word_length*2]};
assign pixels_24_23 = {result[761*word_length*2-1 -: word_length*2]};
assign pixels_25_23 = {result[762*word_length*2-1 -: word_length*2]};
assign pixels_26_23 = {result[763*word_length*2-1 -: word_length*2]};
assign pixels_27_23 = {result[764*word_length*2-1 -: word_length*2]};
assign pixels_28_23 = {result[765*word_length*2-1 -: word_length*2]};
assign pixels_29_23 = {result[766*word_length*2-1 -: word_length*2]};
assign pixels_30_23 = {result[767*word_length*2-1 -: word_length*2]};
assign pixels_31_23 = {result[768*word_length*2-1 -: word_length*2]};
assign pixels_0_24 = {result[769*word_length*2-1 -: word_length*2]};
assign pixels_1_24 = {result[770*word_length*2-1 -: word_length*2]};
assign pixels_2_24 = {result[771*word_length*2-1 -: word_length*2]};
assign pixels_3_24 = {result[772*word_length*2-1 -: word_length*2]};
assign pixels_4_24 = {result[773*word_length*2-1 -: word_length*2]};
assign pixels_5_24 = {result[774*word_length*2-1 -: word_length*2]};
assign pixels_6_24 = {result[775*word_length*2-1 -: word_length*2]};
assign pixels_7_24 = {result[776*word_length*2-1 -: word_length*2]};
assign pixels_8_24 = {result[777*word_length*2-1 -: word_length*2]};
assign pixels_9_24 = {result[778*word_length*2-1 -: word_length*2]};
assign pixels_10_24 = {result[779*word_length*2-1 -: word_length*2]};
assign pixels_11_24 = {result[780*word_length*2-1 -: word_length*2]};
assign pixels_12_24 = {result[781*word_length*2-1 -: word_length*2]};
assign pixels_13_24 = {result[782*word_length*2-1 -: word_length*2]};
assign pixels_14_24 = {result[783*word_length*2-1 -: word_length*2]};
assign pixels_15_24 = {result[784*word_length*2-1 -: word_length*2]};
assign pixels_16_24 = {result[785*word_length*2-1 -: word_length*2]};
assign pixels_17_24 = {result[786*word_length*2-1 -: word_length*2]};
assign pixels_18_24 = {result[787*word_length*2-1 -: word_length*2]};
assign pixels_19_24 = {result[788*word_length*2-1 -: word_length*2]};
assign pixels_20_24 = {result[789*word_length*2-1 -: word_length*2]};
assign pixels_21_24 = {result[790*word_length*2-1 -: word_length*2]};
assign pixels_22_24 = {result[791*word_length*2-1 -: word_length*2]};
assign pixels_23_24 = {result[792*word_length*2-1 -: word_length*2]};
assign pixels_24_24 = {result[793*word_length*2-1 -: word_length*2]};
assign pixels_25_24 = {result[794*word_length*2-1 -: word_length*2]};
assign pixels_26_24 = {result[795*word_length*2-1 -: word_length*2]};
assign pixels_27_24 = {result[796*word_length*2-1 -: word_length*2]};
assign pixels_28_24 = {result[797*word_length*2-1 -: word_length*2]};
assign pixels_29_24 = {result[798*word_length*2-1 -: word_length*2]};
assign pixels_30_24 = {result[799*word_length*2-1 -: word_length*2]};
assign pixels_31_24 = {result[800*word_length*2-1 -: word_length*2]};
assign pixels_0_25 = {result[801*word_length*2-1 -: word_length*2]};
assign pixels_1_25 = {result[802*word_length*2-1 -: word_length*2]};
assign pixels_2_25 = {result[803*word_length*2-1 -: word_length*2]};
assign pixels_3_25 = {result[804*word_length*2-1 -: word_length*2]};
assign pixels_4_25 = {result[805*word_length*2-1 -: word_length*2]};
assign pixels_5_25 = {result[806*word_length*2-1 -: word_length*2]};
assign pixels_6_25 = {result[807*word_length*2-1 -: word_length*2]};
assign pixels_7_25 = {result[808*word_length*2-1 -: word_length*2]};
assign pixels_8_25 = {result[809*word_length*2-1 -: word_length*2]};
assign pixels_9_25 = {result[810*word_length*2-1 -: word_length*2]};
assign pixels_10_25 = {result[811*word_length*2-1 -: word_length*2]};
assign pixels_11_25 = {result[812*word_length*2-1 -: word_length*2]};
assign pixels_12_25 = {result[813*word_length*2-1 -: word_length*2]};
assign pixels_13_25 = {result[814*word_length*2-1 -: word_length*2]};
assign pixels_14_25 = {result[815*word_length*2-1 -: word_length*2]};
assign pixels_15_25 = {result[816*word_length*2-1 -: word_length*2]};
assign pixels_16_25 = {result[817*word_length*2-1 -: word_length*2]};
assign pixels_17_25 = {result[818*word_length*2-1 -: word_length*2]};
assign pixels_18_25 = {result[819*word_length*2-1 -: word_length*2]};
assign pixels_19_25 = {result[820*word_length*2-1 -: word_length*2]};
assign pixels_20_25 = {result[821*word_length*2-1 -: word_length*2]};
assign pixels_21_25 = {result[822*word_length*2-1 -: word_length*2]};
assign pixels_22_25 = {result[823*word_length*2-1 -: word_length*2]};
assign pixels_23_25 = {result[824*word_length*2-1 -: word_length*2]};
assign pixels_24_25 = {result[825*word_length*2-1 -: word_length*2]};
assign pixels_25_25 = {result[826*word_length*2-1 -: word_length*2]};
assign pixels_26_25 = {result[827*word_length*2-1 -: word_length*2]};
assign pixels_27_25 = {result[828*word_length*2-1 -: word_length*2]};
assign pixels_28_25 = {result[829*word_length*2-1 -: word_length*2]};
assign pixels_29_25 = {result[830*word_length*2-1 -: word_length*2]};
assign pixels_30_25 = {result[831*word_length*2-1 -: word_length*2]};
assign pixels_31_25 = {result[832*word_length*2-1 -: word_length*2]};
assign pixels_0_26 = {result[833*word_length*2-1 -: word_length*2]};
assign pixels_1_26 = {result[834*word_length*2-1 -: word_length*2]};
assign pixels_2_26 = {result[835*word_length*2-1 -: word_length*2]};
assign pixels_3_26 = {result[836*word_length*2-1 -: word_length*2]};
assign pixels_4_26 = {result[837*word_length*2-1 -: word_length*2]};
assign pixels_5_26 = {result[838*word_length*2-1 -: word_length*2]};
assign pixels_6_26 = {result[839*word_length*2-1 -: word_length*2]};
assign pixels_7_26 = {result[840*word_length*2-1 -: word_length*2]};
assign pixels_8_26 = {result[841*word_length*2-1 -: word_length*2]};
assign pixels_9_26 = {result[842*word_length*2-1 -: word_length*2]};
assign pixels_10_26 = {result[843*word_length*2-1 -: word_length*2]};
assign pixels_11_26 = {result[844*word_length*2-1 -: word_length*2]};
assign pixels_12_26 = {result[845*word_length*2-1 -: word_length*2]};
assign pixels_13_26 = {result[846*word_length*2-1 -: word_length*2]};
assign pixels_14_26 = {result[847*word_length*2-1 -: word_length*2]};
assign pixels_15_26 = {result[848*word_length*2-1 -: word_length*2]};
assign pixels_16_26 = {result[849*word_length*2-1 -: word_length*2]};
assign pixels_17_26 = {result[850*word_length*2-1 -: word_length*2]};
assign pixels_18_26 = {result[851*word_length*2-1 -: word_length*2]};
assign pixels_19_26 = {result[852*word_length*2-1 -: word_length*2]};
assign pixels_20_26 = {result[853*word_length*2-1 -: word_length*2]};
assign pixels_21_26 = {result[854*word_length*2-1 -: word_length*2]};
assign pixels_22_26 = {result[855*word_length*2-1 -: word_length*2]};
assign pixels_23_26 = {result[856*word_length*2-1 -: word_length*2]};
assign pixels_24_26 = {result[857*word_length*2-1 -: word_length*2]};
assign pixels_25_26 = {result[858*word_length*2-1 -: word_length*2]};
assign pixels_26_26 = {result[859*word_length*2-1 -: word_length*2]};
assign pixels_27_26 = {result[860*word_length*2-1 -: word_length*2]};
assign pixels_28_26 = {result[861*word_length*2-1 -: word_length*2]};
assign pixels_29_26 = {result[862*word_length*2-1 -: word_length*2]};
assign pixels_30_26 = {result[863*word_length*2-1 -: word_length*2]};
assign pixels_31_26 = {result[864*word_length*2-1 -: word_length*2]};
assign pixels_0_27 = {result[865*word_length*2-1 -: word_length*2]};
assign pixels_1_27 = {result[866*word_length*2-1 -: word_length*2]};
assign pixels_2_27 = {result[867*word_length*2-1 -: word_length*2]};
assign pixels_3_27 = {result[868*word_length*2-1 -: word_length*2]};
assign pixels_4_27 = {result[869*word_length*2-1 -: word_length*2]};
assign pixels_5_27 = {result[870*word_length*2-1 -: word_length*2]};
assign pixels_6_27 = {result[871*word_length*2-1 -: word_length*2]};
assign pixels_7_27 = {result[872*word_length*2-1 -: word_length*2]};
assign pixels_8_27 = {result[873*word_length*2-1 -: word_length*2]};
assign pixels_9_27 = {result[874*word_length*2-1 -: word_length*2]};
assign pixels_10_27 = {result[875*word_length*2-1 -: word_length*2]};
assign pixels_11_27 = {result[876*word_length*2-1 -: word_length*2]};
assign pixels_12_27 = {result[877*word_length*2-1 -: word_length*2]};
assign pixels_13_27 = {result[878*word_length*2-1 -: word_length*2]};
assign pixels_14_27 = {result[879*word_length*2-1 -: word_length*2]};
assign pixels_15_27 = {result[880*word_length*2-1 -: word_length*2]};
assign pixels_16_27 = {result[881*word_length*2-1 -: word_length*2]};
assign pixels_17_27 = {result[882*word_length*2-1 -: word_length*2]};
assign pixels_18_27 = {result[883*word_length*2-1 -: word_length*2]};
assign pixels_19_27 = {result[884*word_length*2-1 -: word_length*2]};
assign pixels_20_27 = {result[885*word_length*2-1 -: word_length*2]};
assign pixels_21_27 = {result[886*word_length*2-1 -: word_length*2]};
assign pixels_22_27 = {result[887*word_length*2-1 -: word_length*2]};
assign pixels_23_27 = {result[888*word_length*2-1 -: word_length*2]};
assign pixels_24_27 = {result[889*word_length*2-1 -: word_length*2]};
assign pixels_25_27 = {result[890*word_length*2-1 -: word_length*2]};
assign pixels_26_27 = {result[891*word_length*2-1 -: word_length*2]};
assign pixels_27_27 = {result[892*word_length*2-1 -: word_length*2]};
assign pixels_28_27 = {result[893*word_length*2-1 -: word_length*2]};
assign pixels_29_27 = {result[894*word_length*2-1 -: word_length*2]};
assign pixels_30_27 = {result[895*word_length*2-1 -: word_length*2]};
assign pixels_31_27 = {result[896*word_length*2-1 -: word_length*2]};
assign pixels_0_28 = {result[897*word_length*2-1 -: word_length*2]};
assign pixels_1_28 = {result[898*word_length*2-1 -: word_length*2]};
assign pixels_2_28 = {result[899*word_length*2-1 -: word_length*2]};
assign pixels_3_28 = {result[900*word_length*2-1 -: word_length*2]};
assign pixels_4_28 = {result[901*word_length*2-1 -: word_length*2]};
assign pixels_5_28 = {result[902*word_length*2-1 -: word_length*2]};
assign pixels_6_28 = {result[903*word_length*2-1 -: word_length*2]};
assign pixels_7_28 = {result[904*word_length*2-1 -: word_length*2]};
assign pixels_8_28 = {result[905*word_length*2-1 -: word_length*2]};
assign pixels_9_28 = {result[906*word_length*2-1 -: word_length*2]};
assign pixels_10_28 = {result[907*word_length*2-1 -: word_length*2]};
assign pixels_11_28 = {result[908*word_length*2-1 -: word_length*2]};
assign pixels_12_28 = {result[909*word_length*2-1 -: word_length*2]};
assign pixels_13_28 = {result[910*word_length*2-1 -: word_length*2]};
assign pixels_14_28 = {result[911*word_length*2-1 -: word_length*2]};
assign pixels_15_28 = {result[912*word_length*2-1 -: word_length*2]};
assign pixels_16_28 = {result[913*word_length*2-1 -: word_length*2]};
assign pixels_17_28 = {result[914*word_length*2-1 -: word_length*2]};
assign pixels_18_28 = {result[915*word_length*2-1 -: word_length*2]};
assign pixels_19_28 = {result[916*word_length*2-1 -: word_length*2]};
assign pixels_20_28 = {result[917*word_length*2-1 -: word_length*2]};
assign pixels_21_28 = {result[918*word_length*2-1 -: word_length*2]};
assign pixels_22_28 = {result[919*word_length*2-1 -: word_length*2]};
assign pixels_23_28 = {result[920*word_length*2-1 -: word_length*2]};
assign pixels_24_28 = {result[921*word_length*2-1 -: word_length*2]};
assign pixels_25_28 = {result[922*word_length*2-1 -: word_length*2]};
assign pixels_26_28 = {result[923*word_length*2-1 -: word_length*2]};
assign pixels_27_28 = {result[924*word_length*2-1 -: word_length*2]};
assign pixels_28_28 = {result[925*word_length*2-1 -: word_length*2]};
assign pixels_29_28 = {result[926*word_length*2-1 -: word_length*2]};
assign pixels_30_28 = {result[927*word_length*2-1 -: word_length*2]};
assign pixels_31_28 = {result[928*word_length*2-1 -: word_length*2]};
assign pixels_0_29 = {result[929*word_length*2-1 -: word_length*2]};
assign pixels_1_29 = {result[930*word_length*2-1 -: word_length*2]};
assign pixels_2_29 = {result[931*word_length*2-1 -: word_length*2]};
assign pixels_3_29 = {result[932*word_length*2-1 -: word_length*2]};
assign pixels_4_29 = {result[933*word_length*2-1 -: word_length*2]};
assign pixels_5_29 = {result[934*word_length*2-1 -: word_length*2]};
assign pixels_6_29 = {result[935*word_length*2-1 -: word_length*2]};
assign pixels_7_29 = {result[936*word_length*2-1 -: word_length*2]};
assign pixels_8_29 = {result[937*word_length*2-1 -: word_length*2]};
assign pixels_9_29 = {result[938*word_length*2-1 -: word_length*2]};
assign pixels_10_29 = {result[939*word_length*2-1 -: word_length*2]};
assign pixels_11_29 = {result[940*word_length*2-1 -: word_length*2]};
assign pixels_12_29 = {result[941*word_length*2-1 -: word_length*2]};
assign pixels_13_29 = {result[942*word_length*2-1 -: word_length*2]};
assign pixels_14_29 = {result[943*word_length*2-1 -: word_length*2]};
assign pixels_15_29 = {result[944*word_length*2-1 -: word_length*2]};
assign pixels_16_29 = {result[945*word_length*2-1 -: word_length*2]};
assign pixels_17_29 = {result[946*word_length*2-1 -: word_length*2]};
assign pixels_18_29 = {result[947*word_length*2-1 -: word_length*2]};
assign pixels_19_29 = {result[948*word_length*2-1 -: word_length*2]};
assign pixels_20_29 = {result[949*word_length*2-1 -: word_length*2]};
assign pixels_21_29 = {result[950*word_length*2-1 -: word_length*2]};
assign pixels_22_29 = {result[951*word_length*2-1 -: word_length*2]};
assign pixels_23_29 = {result[952*word_length*2-1 -: word_length*2]};
assign pixels_24_29 = {result[953*word_length*2-1 -: word_length*2]};
assign pixels_25_29 = {result[954*word_length*2-1 -: word_length*2]};
assign pixels_26_29 = {result[955*word_length*2-1 -: word_length*2]};
assign pixels_27_29 = {result[956*word_length*2-1 -: word_length*2]};
assign pixels_28_29 = {result[957*word_length*2-1 -: word_length*2]};
assign pixels_29_29 = {result[958*word_length*2-1 -: word_length*2]};
assign pixels_30_29 = {result[959*word_length*2-1 -: word_length*2]};
assign pixels_31_29 = {result[960*word_length*2-1 -: word_length*2]};
assign pixels_0_30 = {result[961*word_length*2-1 -: word_length*2]};
assign pixels_1_30 = {result[962*word_length*2-1 -: word_length*2]};
assign pixels_2_30 = {result[963*word_length*2-1 -: word_length*2]};
assign pixels_3_30 = {result[964*word_length*2-1 -: word_length*2]};
assign pixels_4_30 = {result[965*word_length*2-1 -: word_length*2]};
assign pixels_5_30 = {result[966*word_length*2-1 -: word_length*2]};
assign pixels_6_30 = {result[967*word_length*2-1 -: word_length*2]};
assign pixels_7_30 = {result[968*word_length*2-1 -: word_length*2]};
assign pixels_8_30 = {result[969*word_length*2-1 -: word_length*2]};
assign pixels_9_30 = {result[970*word_length*2-1 -: word_length*2]};
assign pixels_10_30 = {result[971*word_length*2-1 -: word_length*2]};
assign pixels_11_30 = {result[972*word_length*2-1 -: word_length*2]};
assign pixels_12_30 = {result[973*word_length*2-1 -: word_length*2]};
assign pixels_13_30 = {result[974*word_length*2-1 -: word_length*2]};
assign pixels_14_30 = {result[975*word_length*2-1 -: word_length*2]};
assign pixels_15_30 = {result[976*word_length*2-1 -: word_length*2]};
assign pixels_16_30 = {result[977*word_length*2-1 -: word_length*2]};
assign pixels_17_30 = {result[978*word_length*2-1 -: word_length*2]};
assign pixels_18_30 = {result[979*word_length*2-1 -: word_length*2]};
assign pixels_19_30 = {result[980*word_length*2-1 -: word_length*2]};
assign pixels_20_30 = {result[981*word_length*2-1 -: word_length*2]};
assign pixels_21_30 = {result[982*word_length*2-1 -: word_length*2]};
assign pixels_22_30 = {result[983*word_length*2-1 -: word_length*2]};
assign pixels_23_30 = {result[984*word_length*2-1 -: word_length*2]};
assign pixels_24_30 = {result[985*word_length*2-1 -: word_length*2]};
assign pixels_25_30 = {result[986*word_length*2-1 -: word_length*2]};
assign pixels_26_30 = {result[987*word_length*2-1 -: word_length*2]};
assign pixels_27_30 = {result[988*word_length*2-1 -: word_length*2]};
assign pixels_28_30 = {result[989*word_length*2-1 -: word_length*2]};
assign pixels_29_30 = {result[990*word_length*2-1 -: word_length*2]};
assign pixels_30_30 = {result[991*word_length*2-1 -: word_length*2]};
assign pixels_31_30 = {result[992*word_length*2-1 -: word_length*2]};
assign pixels_0_31 = {result[993*word_length*2-1 -: word_length*2]};
assign pixels_1_31 = {result[994*word_length*2-1 -: word_length*2]};
assign pixels_2_31 = {result[995*word_length*2-1 -: word_length*2]};
assign pixels_3_31 = {result[996*word_length*2-1 -: word_length*2]};
assign pixels_4_31 = {result[997*word_length*2-1 -: word_length*2]};
assign pixels_5_31 = {result[998*word_length*2-1 -: word_length*2]};
assign pixels_6_31 = {result[999*word_length*2-1 -: word_length*2]};
assign pixels_7_31 = {result[1000*word_length*2-1 -: word_length*2]};
assign pixels_8_31 = {result[1001*word_length*2-1 -: word_length*2]};
assign pixels_9_31 = {result[1002*word_length*2-1 -: word_length*2]};
assign pixels_10_31 = {result[1003*word_length*2-1 -: word_length*2]};
assign pixels_11_31 = {result[1004*word_length*2-1 -: word_length*2]};
assign pixels_12_31 = {result[1005*word_length*2-1 -: word_length*2]};
assign pixels_13_31 = {result[1006*word_length*2-1 -: word_length*2]};
assign pixels_14_31 = {result[1007*word_length*2-1 -: word_length*2]};
assign pixels_15_31 = {result[1008*word_length*2-1 -: word_length*2]};
assign pixels_16_31 = {result[1009*word_length*2-1 -: word_length*2]};
assign pixels_17_31 = {result[1010*word_length*2-1 -: word_length*2]};
assign pixels_18_31 = {result[1011*word_length*2-1 -: word_length*2]};
assign pixels_19_31 = {result[1012*word_length*2-1 -: word_length*2]};
assign pixels_20_31 = {result[1013*word_length*2-1 -: word_length*2]};
assign pixels_21_31 = {result[1014*word_length*2-1 -: word_length*2]};
assign pixels_22_31 = {result[1015*word_length*2-1 -: word_length*2]};
assign pixels_23_31 = {result[1016*word_length*2-1 -: word_length*2]};
assign pixels_24_31 = {result[1017*word_length*2-1 -: word_length*2]};
assign pixels_25_31 = {result[1018*word_length*2-1 -: word_length*2]};
assign pixels_26_31 = {result[1019*word_length*2-1 -: word_length*2]};
assign pixels_27_31 = {result[1020*word_length*2-1 -: word_length*2]};
assign pixels_28_31 = {result[1021*word_length*2-1 -: word_length*2]};
assign pixels_29_31 = {result[1022*word_length*2-1 -: word_length*2]};
assign pixels_30_31 = {result[1023*word_length*2-1 -: word_length*2]};
assign pixels_31_31 = {result[1024*word_length*2-1 -: word_length*2]};

//iter
integer i,j;

initial begin
    #0      rst = 0;
            clk = 1;
            feature_valid_num = 16'd195;
            weight_valid_num = 16'd27;
            result = 0;
            $display("START!\n");
    #10     rst = 1;
    #10     rst = 0;
    #100    in_valid = 1;

    #16000  
if(pixels_0_0!==16'hffb6) $display("ERROR! at (0,0)\n");
if(pixels_1_0!==16'hfd25) $display("ERROR! at (1,0)\n");
if(pixels_2_0!==16'hfd93) $display("ERROR! at (2,0)\n");
if(pixels_3_0!==16'hfed3) $display("ERROR! at (3,0)\n");
if(pixels_4_0!==16'h0337) $display("ERROR! at (4,0)\n");
if(pixels_5_0!==16'h02ba) $display("ERROR! at (5,0)\n");
if(pixels_6_0!==16'hfde6) $display("ERROR! at (6,0)\n");
if(pixels_7_0!==16'h00d0) $display("ERROR! at (7,0)\n");
if(pixels_8_0!==16'h01a7) $display("ERROR! at (8,0)\n");
if(pixels_9_0!==16'h088e) $display("ERROR! at (9,0)\n");
if(pixels_10_0!==16'h01ed) $display("ERROR! at (10,0)\n");
if(pixels_11_0!==16'h0365) $display("ERROR! at (11,0)\n");
if(pixels_12_0!==16'hfb29) $display("ERROR! at (12,0)\n");
if(pixels_13_0!==16'h011c) $display("ERROR! at (13,0)\n");
if(pixels_14_0!==16'hff2e) $display("ERROR! at (14,0)\n");
if(pixels_15_0!==16'h0139) $display("ERROR! at (15,0)\n");
if(pixels_16_0!==16'hfd31) $display("ERROR! at (16,0)\n");
if(pixels_17_0!==16'hffe3) $display("ERROR! at (17,0)\n");
if(pixels_18_0!==16'h00ef) $display("ERROR! at (18,0)\n");
if(pixels_19_0!==16'h0032) $display("ERROR! at (19,0)\n");
if(pixels_20_0!==16'h029e) $display("ERROR! at (20,0)\n");
if(pixels_21_0!==16'hffd6) $display("ERROR! at (21,0)\n");
if(pixels_22_0!==16'h00db) $display("ERROR! at (22,0)\n");
if(pixels_23_0!==16'h02fb) $display("ERROR! at (23,0)\n");
if(pixels_24_0!==16'h0124) $display("ERROR! at (24,0)\n");
if(pixels_25_0!==16'hfe0d) $display("ERROR! at (25,0)\n");
if(pixels_26_0!==16'hfd3c) $display("ERROR! at (26,0)\n");
if(pixels_27_0!==16'h02ab) $display("ERROR! at (27,0)\n");
if(pixels_28_0!==16'h00c1) $display("ERROR! at (28,0)\n");
if(pixels_29_0!==16'hffde) $display("ERROR! at (29,0)\n");
if(pixels_30_0!==16'hff29) $display("ERROR! at (30,0)\n");
if(pixels_31_0!==16'h0096) $display("ERROR! at (31,0)\n");
if(pixels_0_1!==16'hfe3c) $display("ERROR! at (0,1)\n");
if(pixels_1_1!==16'hfeed) $display("ERROR! at (1,1)\n");
if(pixels_2_1!==16'hff52) $display("ERROR! at (2,1)\n");
if(pixels_3_1!==16'h057e) $display("ERROR! at (3,1)\n");
if(pixels_4_1!==16'hfd70) $display("ERROR! at (4,1)\n");
if(pixels_5_1!==16'hfe18) $display("ERROR! at (5,1)\n");
if(pixels_6_1!==16'hf527) $display("ERROR! at (6,1)\n");
if(pixels_7_1!==16'h006f) $display("ERROR! at (7,1)\n");
if(pixels_8_1!==16'h0300) $display("ERROR! at (8,1)\n");
if(pixels_9_1!==16'hfd6c) $display("ERROR! at (9,1)\n");
if(pixels_10_1!==16'h00fa) $display("ERROR! at (10,1)\n");
if(pixels_11_1!==16'hf60d) $display("ERROR! at (11,1)\n");
if(pixels_12_1!==16'hf50f) $display("ERROR! at (12,1)\n");
if(pixels_13_1!==16'hffaf) $display("ERROR! at (13,1)\n");
if(pixels_14_1!==16'h00f5) $display("ERROR! at (14,1)\n");
if(pixels_15_1!==16'h009b) $display("ERROR! at (15,1)\n");
if(pixels_16_1!==16'h0039) $display("ERROR! at (16,1)\n");
if(pixels_17_1!==16'hff85) $display("ERROR! at (17,1)\n");
if(pixels_18_1!==16'h00a7) $display("ERROR! at (18,1)\n");
if(pixels_19_1!==16'h0454) $display("ERROR! at (19,1)\n");
if(pixels_20_1!==16'hfe3a) $display("ERROR! at (20,1)\n");
if(pixels_21_1!==16'hf85e) $display("ERROR! at (21,1)\n");
if(pixels_22_1!==16'hfc58) $display("ERROR! at (22,1)\n");
if(pixels_23_1!==16'h001f) $display("ERROR! at (23,1)\n");
if(pixels_24_1!==16'hf88c) $display("ERROR! at (24,1)\n");
if(pixels_25_1!==16'hfaa1) $display("ERROR! at (25,1)\n");
if(pixels_26_1!==16'h0071) $display("ERROR! at (26,1)\n");
if(pixels_27_1!==16'h0210) $display("ERROR! at (27,1)\n");
if(pixels_28_1!==16'hfef0) $display("ERROR! at (28,1)\n");
if(pixels_29_1!==16'hffe3) $display("ERROR! at (29,1)\n");
if(pixels_30_1!==16'hffa4) $display("ERROR! at (30,1)\n");
if(pixels_31_1!==16'hffab) $display("ERROR! at (31,1)\n");
if(pixels_0_2!==16'hfae8) $display("ERROR! at (0,2)\n");
if(pixels_1_2!==16'h0267) $display("ERROR! at (1,2)\n");
if(pixels_2_2!==16'hffe2) $display("ERROR! at (2,2)\n");
if(pixels_3_2!==16'h06d0) $display("ERROR! at (3,2)\n");
if(pixels_4_2!==16'hf9d9) $display("ERROR! at (4,2)\n");
if(pixels_5_2!==16'hfb86) $display("ERROR! at (5,2)\n");
if(pixels_6_2!==16'h0226) $display("ERROR! at (6,2)\n");
if(pixels_7_2!==16'h047e) $display("ERROR! at (7,2)\n");
if(pixels_8_2!==16'hfe12) $display("ERROR! at (8,2)\n");
if(pixels_9_2!==16'h069b) $display("ERROR! at (9,2)\n");
if(pixels_10_2!==16'hf6b5) $display("ERROR! at (10,2)\n");
if(pixels_11_2!==16'h04ea) $display("ERROR! at (11,2)\n");
if(pixels_12_2!==16'hf66c) $display("ERROR! at (12,2)\n");
if(pixels_13_2!==16'h05e2) $display("ERROR! at (13,2)\n");
if(pixels_14_2!==16'hfe7e) $display("ERROR! at (14,2)\n");
if(pixels_15_2!==16'h0bfd) $display("ERROR! at (15,2)\n");
if(pixels_16_2!==16'hfbd9) $display("ERROR! at (16,2)\n");
if(pixels_17_2!==16'hfc46) $display("ERROR! at (17,2)\n");
if(pixels_18_2!==16'h033b) $display("ERROR! at (18,2)\n");
if(pixels_19_2!==16'hfb2c) $display("ERROR! at (19,2)\n");
if(pixels_20_2!==16'hfce7) $display("ERROR! at (20,2)\n");
if(pixels_21_2!==16'hf98b) $display("ERROR! at (21,2)\n");
if(pixels_22_2!==16'h0131) $display("ERROR! at (22,2)\n");
if(pixels_23_2!==16'hfecd) $display("ERROR! at (23,2)\n");
if(pixels_24_2!==16'h063f) $display("ERROR! at (24,2)\n");
if(pixels_25_2!==16'h0901) $display("ERROR! at (25,2)\n");
if(pixels_26_2!==16'h0290) $display("ERROR! at (26,2)\n");
if(pixels_27_2!==16'hfb6d) $display("ERROR! at (27,2)\n");
if(pixels_28_2!==16'hff8e) $display("ERROR! at (28,2)\n");
if(pixels_29_2!==16'h016f) $display("ERROR! at (29,2)\n");
if(pixels_30_2!==16'h01ea) $display("ERROR! at (30,2)\n");
if(pixels_31_2!==16'hfd95) $display("ERROR! at (31,2)\n");
if(pixels_0_3!==16'hfdab) $display("ERROR! at (0,3)\n");
if(pixels_1_3!==16'h05f7) $display("ERROR! at (1,3)\n");
if(pixels_2_3!==16'h06c2) $display("ERROR! at (2,3)\n");
if(pixels_3_3!==16'h02d4) $display("ERROR! at (3,3)\n");
if(pixels_4_3!==16'hee27) $display("ERROR! at (4,3)\n");
if(pixels_5_3!==16'hff0b) $display("ERROR! at (5,3)\n");
if(pixels_6_3!==16'hfef3) $display("ERROR! at (6,3)\n");
if(pixels_7_3!==16'h07e4) $display("ERROR! at (7,3)\n");
if(pixels_8_3!==16'hfd7c) $display("ERROR! at (8,3)\n");
if(pixels_9_3!==16'hf72b) $display("ERROR! at (9,3)\n");
if(pixels_10_3!==16'h078f) $display("ERROR! at (10,3)\n");
if(pixels_11_3!==16'h05b4) $display("ERROR! at (11,3)\n");
if(pixels_12_3!==16'hfed1) $display("ERROR! at (12,3)\n");
if(pixels_13_3!==16'h013d) $display("ERROR! at (13,3)\n");
if(pixels_14_3!==16'hf684) $display("ERROR! at (14,3)\n");
if(pixels_15_3!==16'hfed8) $display("ERROR! at (15,3)\n");
if(pixels_16_3!==16'hf9a8) $display("ERROR! at (16,3)\n");
if(pixels_17_3!==16'hfa8b) $display("ERROR! at (17,3)\n");
if(pixels_18_3!==16'hfe86) $display("ERROR! at (18,3)\n");
if(pixels_19_3!==16'hfd03) $display("ERROR! at (19,3)\n");
if(pixels_20_3!==16'h039c) $display("ERROR! at (20,3)\n");
if(pixels_21_3!==16'hfe82) $display("ERROR! at (21,3)\n");
if(pixels_22_3!==16'h0452) $display("ERROR! at (22,3)\n");
if(pixels_23_3!==16'h048e) $display("ERROR! at (23,3)\n");
if(pixels_24_3!==16'h0a41) $display("ERROR! at (24,3)\n");
if(pixels_25_3!==16'h07df) $display("ERROR! at (25,3)\n");
if(pixels_26_3!==16'hfa4d) $display("ERROR! at (26,3)\n");
if(pixels_27_3!==16'hfa2e) $display("ERROR! at (27,3)\n");
if(pixels_28_3!==16'h03c3) $display("ERROR! at (28,3)\n");
if(pixels_29_3!==16'h03ad) $display("ERROR! at (29,3)\n");
if(pixels_30_3!==16'hffda) $display("ERROR! at (30,3)\n");
if(pixels_31_3!==16'h027c) $display("ERROR! at (31,3)\n");
if(pixels_0_4!==16'h01bd) $display("ERROR! at (0,4)\n");
if(pixels_1_4!==16'hff72) $display("ERROR! at (1,4)\n");
if(pixels_2_4!==16'hfd11) $display("ERROR! at (2,4)\n");
if(pixels_3_4!==16'hfd93) $display("ERROR! at (3,4)\n");
if(pixels_4_4!==16'hfdc0) $display("ERROR! at (4,4)\n");
if(pixels_5_4!==16'h0300) $display("ERROR! at (5,4)\n");
if(pixels_6_4!==16'h02b0) $display("ERROR! at (6,4)\n");
if(pixels_7_4!==16'hfc42) $display("ERROR! at (7,4)\n");
if(pixels_8_4!==16'hfc19) $display("ERROR! at (8,4)\n");
if(pixels_9_4!==16'hff57) $display("ERROR! at (9,4)\n");
if(pixels_10_4!==16'h05bb) $display("ERROR! at (10,4)\n");
if(pixels_11_4!==16'h0266) $display("ERROR! at (11,4)\n");
if(pixels_12_4!==16'hfc67) $display("ERROR! at (12,4)\n");
if(pixels_13_4!==16'hfefc) $display("ERROR! at (13,4)\n");
if(pixels_14_4!==16'hf91d) $display("ERROR! at (14,4)\n");
if(pixels_15_4!==16'hff5f) $display("ERROR! at (15,4)\n");
if(pixels_16_4!==16'h0e65) $display("ERROR! at (16,4)\n");
if(pixels_17_4!==16'h035c) $display("ERROR! at (17,4)\n");
if(pixels_18_4!==16'h058f) $display("ERROR! at (18,4)\n");
if(pixels_19_4!==16'h046c) $display("ERROR! at (19,4)\n");
if(pixels_20_4!==16'h09fb) $display("ERROR! at (20,4)\n");
if(pixels_21_4!==16'h01b4) $display("ERROR! at (21,4)\n");
if(pixels_22_4!==16'h02f0) $display("ERROR! at (22,4)\n");
if(pixels_23_4!==16'h0298) $display("ERROR! at (23,4)\n");
if(pixels_24_4!==16'h0103) $display("ERROR! at (24,4)\n");
if(pixels_25_4!==16'hfd33) $display("ERROR! at (25,4)\n");
if(pixels_26_4!==16'hfd4d) $display("ERROR! at (26,4)\n");
if(pixels_27_4!==16'hf89d) $display("ERROR! at (27,4)\n");
if(pixels_28_4!==16'hf552) $display("ERROR! at (28,4)\n");
if(pixels_29_4!==16'hfc0c) $display("ERROR! at (29,4)\n");
if(pixels_30_4!==16'h05b8) $display("ERROR! at (30,4)\n");
if(pixels_31_4!==16'hfc77) $display("ERROR! at (31,4)\n");
if(pixels_0_5!==16'hfe2a) $display("ERROR! at (0,5)\n");
if(pixels_1_5!==16'hfb4a) $display("ERROR! at (1,5)\n");
if(pixels_2_5!==16'h002b) $display("ERROR! at (2,5)\n");
if(pixels_3_5!==16'h04be) $display("ERROR! at (3,5)\n");
if(pixels_4_5!==16'h061a) $display("ERROR! at (4,5)\n");
if(pixels_5_5!==16'h04fc) $display("ERROR! at (5,5)\n");
if(pixels_6_5!==16'h0338) $display("ERROR! at (6,5)\n");
if(pixels_7_5!==16'h027b) $display("ERROR! at (7,5)\n");
if(pixels_8_5!==16'hfe34) $display("ERROR! at (8,5)\n");
if(pixels_9_5!==16'hfc12) $display("ERROR! at (9,5)\n");
if(pixels_10_5!==16'h017c) $display("ERROR! at (10,5)\n");
if(pixels_11_5!==16'hffbc) $display("ERROR! at (11,5)\n");
if(pixels_12_5!==16'hfe6d) $display("ERROR! at (12,5)\n");
if(pixels_13_5!==16'h0502) $display("ERROR! at (13,5)\n");
if(pixels_14_5!==16'hfdc3) $display("ERROR! at (14,5)\n");
if(pixels_15_5!==16'h0d15) $display("ERROR! at (15,5)\n");
if(pixels_16_5!==16'h06a3) $display("ERROR! at (16,5)\n");
if(pixels_17_5!==16'h01da) $display("ERROR! at (17,5)\n");
if(pixels_18_5!==16'h0307) $display("ERROR! at (18,5)\n");
if(pixels_19_5!==16'h03a3) $display("ERROR! at (19,5)\n");
if(pixels_20_5!==16'h0155) $display("ERROR! at (20,5)\n");
if(pixels_21_5!==16'hf30b) $display("ERROR! at (21,5)\n");
if(pixels_22_5!==16'hf9b8) $display("ERROR! at (22,5)\n");
if(pixels_23_5!==16'hfd18) $display("ERROR! at (23,5)\n");
if(pixels_24_5!==16'h007b) $display("ERROR! at (24,5)\n");
if(pixels_25_5!==16'h03dd) $display("ERROR! at (25,5)\n");
if(pixels_26_5!==16'h035f) $display("ERROR! at (26,5)\n");
if(pixels_27_5!==16'hf61a) $display("ERROR! at (27,5)\n");
if(pixels_28_5!==16'h0b15) $display("ERROR! at (28,5)\n");
if(pixels_29_5!==16'h045c) $display("ERROR! at (29,5)\n");
if(pixels_30_5!==16'hfcc5) $display("ERROR! at (30,5)\n");
if(pixels_31_5!==16'h0200) $display("ERROR! at (31,5)\n");
if(pixels_0_6!==16'hfcc5) $display("ERROR! at (0,6)\n");
if(pixels_1_6!==16'h0392) $display("ERROR! at (1,6)\n");
if(pixels_2_6!==16'h01c6) $display("ERROR! at (2,6)\n");
if(pixels_3_6!==16'hfe2c) $display("ERROR! at (3,6)\n");
if(pixels_4_6!==16'h005b) $display("ERROR! at (4,6)\n");
if(pixels_5_6!==16'hfe6c) $display("ERROR! at (5,6)\n");
if(pixels_6_6!==16'h0035) $display("ERROR! at (6,6)\n");
if(pixels_7_6!==16'hf88d) $display("ERROR! at (7,6)\n");
if(pixels_8_6!==16'hfec6) $display("ERROR! at (8,6)\n");
if(pixels_9_6!==16'hfe38) $display("ERROR! at (9,6)\n");
if(pixels_10_6!==16'hfa32) $display("ERROR! at (10,6)\n");
if(pixels_11_6!==16'hfea1) $display("ERROR! at (11,6)\n");
if(pixels_12_6!==16'hff12) $display("ERROR! at (12,6)\n");
if(pixels_13_6!==16'hfdb2) $display("ERROR! at (13,6)\n");
if(pixels_14_6!==16'hfdd5) $display("ERROR! at (14,6)\n");
if(pixels_15_6!==16'h011f) $display("ERROR! at (15,6)\n");
if(pixels_16_6!==16'hf672) $display("ERROR! at (16,6)\n");
if(pixels_17_6!==16'hf511) $display("ERROR! at (17,6)\n");
if(pixels_18_6!==16'h0613) $display("ERROR! at (18,6)\n");
if(pixels_19_6!==16'hf825) $display("ERROR! at (19,6)\n");
if(pixels_20_6!==16'hfdc9) $display("ERROR! at (20,6)\n");
if(pixels_21_6!==16'hfc0f) $display("ERROR! at (21,6)\n");
if(pixels_22_6!==16'hffb2) $display("ERROR! at (22,6)\n");
if(pixels_23_6!==16'hfd7a) $display("ERROR! at (23,6)\n");
if(pixels_24_6!==16'h0265) $display("ERROR! at (24,6)\n");
if(pixels_25_6!==16'h075c) $display("ERROR! at (25,6)\n");
if(pixels_26_6!==16'hfe34) $display("ERROR! at (26,6)\n");
if(pixels_27_6!==16'hff04) $display("ERROR! at (27,6)\n");
if(pixels_28_6!==16'hf974) $display("ERROR! at (28,6)\n");
if(pixels_29_6!==16'hf845) $display("ERROR! at (29,6)\n");
if(pixels_30_6!==16'h0717) $display("ERROR! at (30,6)\n");
if(pixels_31_6!==16'h02ef) $display("ERROR! at (31,6)\n");
if(pixels_0_7!==16'hfa71) $display("ERROR! at (0,7)\n");
if(pixels_1_7!==16'h0418) $display("ERROR! at (1,7)\n");
if(pixels_2_7!==16'hfdaf) $display("ERROR! at (2,7)\n");
if(pixels_3_7!==16'hfc3a) $display("ERROR! at (3,7)\n");
if(pixels_4_7!==16'h04a1) $display("ERROR! at (4,7)\n");
if(pixels_5_7!==16'h07b4) $display("ERROR! at (5,7)\n");
if(pixels_6_7!==16'hff25) $display("ERROR! at (6,7)\n");
if(pixels_7_7!==16'h0168) $display("ERROR! at (7,7)\n");
if(pixels_8_7!==16'h03cc) $display("ERROR! at (8,7)\n");
if(pixels_9_7!==16'h05c4) $display("ERROR! at (9,7)\n");
if(pixels_10_7!==16'hffde) $display("ERROR! at (10,7)\n");
if(pixels_11_7!==16'hfebe) $display("ERROR! at (11,7)\n");
if(pixels_12_7!==16'h08e2) $display("ERROR! at (12,7)\n");
if(pixels_13_7!==16'hfb3f) $display("ERROR! at (13,7)\n");
if(pixels_14_7!==16'hf78e) $display("ERROR! at (14,7)\n");
if(pixels_15_7!==16'h033c) $display("ERROR! at (15,7)\n");
if(pixels_16_7!==16'h0cba) $display("ERROR! at (16,7)\n");
if(pixels_17_7!==16'h0aa2) $display("ERROR! at (17,7)\n");
if(pixels_18_7!==16'h0404) $display("ERROR! at (18,7)\n");
if(pixels_19_7!==16'hff3d) $display("ERROR! at (19,7)\n");
if(pixels_20_7!==16'h0219) $display("ERROR! at (20,7)\n");
if(pixels_21_7!==16'h044f) $display("ERROR! at (21,7)\n");
if(pixels_22_7!==16'h0959) $display("ERROR! at (22,7)\n");
if(pixels_23_7!==16'h0131) $display("ERROR! at (23,7)\n");
if(pixels_24_7!==16'h03c3) $display("ERROR! at (24,7)\n");
if(pixels_25_7!==16'h0341) $display("ERROR! at (25,7)\n");
if(pixels_26_7!==16'h035f) $display("ERROR! at (26,7)\n");
if(pixels_27_7!==16'hfa5e) $display("ERROR! at (27,7)\n");
if(pixels_28_7!==16'h0045) $display("ERROR! at (28,7)\n");
if(pixels_29_7!==16'hfdf7) $display("ERROR! at (29,7)\n");
if(pixels_30_7!==16'hf945) $display("ERROR! at (30,7)\n");
if(pixels_31_7!==16'hff7f) $display("ERROR! at (31,7)\n");
if(pixels_0_8!==16'hfcae) $display("ERROR! at (0,8)\n");
if(pixels_1_8!==16'h0632) $display("ERROR! at (1,8)\n");
if(pixels_2_8!==16'h0334) $display("ERROR! at (2,8)\n");
if(pixels_3_8!==16'hfec7) $display("ERROR! at (3,8)\n");
if(pixels_4_8!==16'h0787) $display("ERROR! at (4,8)\n");
if(pixels_5_8!==16'hffbc) $display("ERROR! at (5,8)\n");
if(pixels_6_8!==16'hfe4b) $display("ERROR! at (6,8)\n");
if(pixels_7_8!==16'h064b) $display("ERROR! at (7,8)\n");
if(pixels_8_8!==16'h0661) $display("ERROR! at (8,8)\n");
if(pixels_9_8!==16'h0201) $display("ERROR! at (9,8)\n");
if(pixels_10_8!==16'hfcdd) $display("ERROR! at (10,8)\n");
if(pixels_11_8!==16'h01a4) $display("ERROR! at (11,8)\n");
if(pixels_12_8!==16'hf751) $display("ERROR! at (12,8)\n");
if(pixels_13_8!==16'hf757) $display("ERROR! at (13,8)\n");
if(pixels_14_8!==16'hfcbc) $display("ERROR! at (14,8)\n");
if(pixels_15_8!==16'h044e) $display("ERROR! at (15,8)\n");
if(pixels_16_8!==16'h0b63) $display("ERROR! at (16,8)\n");
if(pixels_17_8!==16'h06e3) $display("ERROR! at (17,8)\n");
if(pixels_18_8!==16'h02fa) $display("ERROR! at (18,8)\n");
if(pixels_19_8!==16'hf4b9) $display("ERROR! at (19,8)\n");
if(pixels_20_8!==16'hf873) $display("ERROR! at (20,8)\n");
if(pixels_21_8!==16'h068e) $display("ERROR! at (21,8)\n");
if(pixels_22_8!==16'hfd0e) $display("ERROR! at (22,8)\n");
if(pixels_23_8!==16'h024a) $display("ERROR! at (23,8)\n");
if(pixels_24_8!==16'hf893) $display("ERROR! at (24,8)\n");
if(pixels_25_8!==16'hfe5f) $display("ERROR! at (25,8)\n");
if(pixels_26_8!==16'hff95) $display("ERROR! at (26,8)\n");
if(pixels_27_8!==16'h0b1c) $display("ERROR! at (27,8)\n");
if(pixels_28_8!==16'h02ad) $display("ERROR! at (28,8)\n");
if(pixels_29_8!==16'hfe6b) $display("ERROR! at (29,8)\n");
if(pixels_30_8!==16'h0166) $display("ERROR! at (30,8)\n");
if(pixels_31_8!==16'h0684) $display("ERROR! at (31,8)\n");
if(pixels_0_9!==16'h010a) $display("ERROR! at (0,9)\n");
if(pixels_1_9!==16'hfb6f) $display("ERROR! at (1,9)\n");
if(pixels_2_9!==16'hfad9) $display("ERROR! at (2,9)\n");
if(pixels_3_9!==16'h061b) $display("ERROR! at (3,9)\n");
if(pixels_4_9!==16'hfb3d) $display("ERROR! at (4,9)\n");
if(pixels_5_9!==16'hf0ba) $display("ERROR! at (5,9)\n");
if(pixels_6_9!==16'h010a) $display("ERROR! at (6,9)\n");
if(pixels_7_9!==16'hfc04) $display("ERROR! at (7,9)\n");
if(pixels_8_9!==16'hfded) $display("ERROR! at (8,9)\n");
if(pixels_9_9!==16'hfd5c) $display("ERROR! at (9,9)\n");
if(pixels_10_9!==16'h03fb) $display("ERROR! at (10,9)\n");
if(pixels_11_9!==16'hf909) $display("ERROR! at (11,9)\n");
if(pixels_12_9!==16'hfdcb) $display("ERROR! at (12,9)\n");
if(pixels_13_9!==16'h0576) $display("ERROR! at (13,9)\n");
if(pixels_14_9!==16'h01e5) $display("ERROR! at (14,9)\n");
if(pixels_15_9!==16'h0031) $display("ERROR! at (15,9)\n");
if(pixels_16_9!==16'hf951) $display("ERROR! at (16,9)\n");
if(pixels_17_9!==16'h0c92) $display("ERROR! at (17,9)\n");
if(pixels_18_9!==16'h0143) $display("ERROR! at (18,9)\n");
if(pixels_19_9!==16'hfc08) $display("ERROR! at (19,9)\n");
if(pixels_20_9!==16'h02e3) $display("ERROR! at (20,9)\n");
if(pixels_21_9!==16'hfda0) $display("ERROR! at (21,9)\n");
if(pixels_22_9!==16'h00e1) $display("ERROR! at (22,9)\n");
if(pixels_23_9!==16'h00da) $display("ERROR! at (23,9)\n");
if(pixels_24_9!==16'hfa5b) $display("ERROR! at (24,9)\n");
if(pixels_25_9!==16'h0559) $display("ERROR! at (25,9)\n");
if(pixels_26_9!==16'h0649) $display("ERROR! at (26,9)\n");
if(pixels_27_9!==16'hfd82) $display("ERROR! at (27,9)\n");
if(pixels_28_9!==16'hfd82) $display("ERROR! at (28,9)\n");
if(pixels_29_9!==16'hf91e) $display("ERROR! at (29,9)\n");
if(pixels_30_9!==16'hff49) $display("ERROR! at (30,9)\n");
if(pixels_31_9!==16'hfe69) $display("ERROR! at (31,9)\n");
if(pixels_0_10!==16'h0415) $display("ERROR! at (0,10)\n");
if(pixels_1_10!==16'hf8bf) $display("ERROR! at (1,10)\n");
if(pixels_2_10!==16'h00e1) $display("ERROR! at (2,10)\n");
if(pixels_3_10!==16'hffe2) $display("ERROR! at (3,10)\n");
if(pixels_4_10!==16'hfdc9) $display("ERROR! at (4,10)\n");
if(pixels_5_10!==16'h0755) $display("ERROR! at (5,10)\n");
if(pixels_6_10!==16'h0530) $display("ERROR! at (6,10)\n");
if(pixels_7_10!==16'hfdc8) $display("ERROR! at (7,10)\n");
if(pixels_8_10!==16'hff36) $display("ERROR! at (8,10)\n");
if(pixels_9_10!==16'hffbf) $display("ERROR! at (9,10)\n");
if(pixels_10_10!==16'hfeb3) $display("ERROR! at (10,10)\n");
if(pixels_11_10!==16'hfea0) $display("ERROR! at (11,10)\n");
if(pixels_12_10!==16'h03ea) $display("ERROR! at (12,10)\n");
if(pixels_13_10!==16'h0beb) $display("ERROR! at (13,10)\n");
if(pixels_14_10!==16'hfb3e) $display("ERROR! at (14,10)\n");
if(pixels_15_10!==16'h0039) $display("ERROR! at (15,10)\n");
if(pixels_16_10!==16'hfec6) $display("ERROR! at (16,10)\n");
if(pixels_17_10!==16'h04ed) $display("ERROR! at (17,10)\n");
if(pixels_18_10!==16'h08a3) $display("ERROR! at (18,10)\n");
if(pixels_19_10!==16'h08a3) $display("ERROR! at (19,10)\n");
if(pixels_20_10!==16'h0102) $display("ERROR! at (20,10)\n");
if(pixels_21_10!==16'hf919) $display("ERROR! at (21,10)\n");
if(pixels_22_10!==16'h0186) $display("ERROR! at (22,10)\n");
if(pixels_23_10!==16'hfea2) $display("ERROR! at (23,10)\n");
if(pixels_24_10!==16'hfebd) $display("ERROR! at (24,10)\n");
if(pixels_25_10!==16'h0840) $display("ERROR! at (25,10)\n");
if(pixels_26_10!==16'hfc96) $display("ERROR! at (26,10)\n");
if(pixels_27_10!==16'h07e7) $display("ERROR! at (27,10)\n");
if(pixels_28_10!==16'hfdbd) $display("ERROR! at (28,10)\n");
if(pixels_29_10!==16'hfe3e) $display("ERROR! at (29,10)\n");
if(pixels_30_10!==16'hfb49) $display("ERROR! at (30,10)\n");
if(pixels_31_10!==16'h0319) $display("ERROR! at (31,10)\n");
if(pixels_0_11!==16'h01b8) $display("ERROR! at (0,11)\n");
if(pixels_1_11!==16'hf91e) $display("ERROR! at (1,11)\n");
if(pixels_2_11!==16'hfc73) $display("ERROR! at (2,11)\n");
if(pixels_3_11!==16'hff57) $display("ERROR! at (3,11)\n");
if(pixels_4_11!==16'hfc38) $display("ERROR! at (4,11)\n");
if(pixels_5_11!==16'h09de) $display("ERROR! at (5,11)\n");
if(pixels_6_11!==16'h074a) $display("ERROR! at (6,11)\n");
if(pixels_7_11!==16'h01d0) $display("ERROR! at (7,11)\n");
if(pixels_8_11!==16'h02bd) $display("ERROR! at (8,11)\n");
if(pixels_9_11!==16'hfd83) $display("ERROR! at (9,11)\n");
if(pixels_10_11!==16'hf9c2) $display("ERROR! at (10,11)\n");
if(pixels_11_11!==16'hfebc) $display("ERROR! at (11,11)\n");
if(pixels_12_11!==16'h0284) $display("ERROR! at (12,11)\n");
if(pixels_13_11!==16'h00ca) $display("ERROR! at (13,11)\n");
if(pixels_14_11!==16'hf788) $display("ERROR! at (14,11)\n");
if(pixels_15_11!==16'h05f8) $display("ERROR! at (15,11)\n");
if(pixels_16_11!==16'hf36e) $display("ERROR! at (16,11)\n");
if(pixels_17_11!==16'h081d) $display("ERROR! at (17,11)\n");
if(pixels_18_11!==16'h0c26) $display("ERROR! at (18,11)\n");
if(pixels_19_11!==16'hf9ff) $display("ERROR! at (19,11)\n");
if(pixels_20_11!==16'hf9ff) $display("ERROR! at (20,11)\n");
if(pixels_21_11!==16'h0181) $display("ERROR! at (21,11)\n");
if(pixels_22_11!==16'hf722) $display("ERROR! at (22,11)\n");
if(pixels_23_11!==16'h0323) $display("ERROR! at (23,11)\n");
if(pixels_24_11!==16'hf6cd) $display("ERROR! at (24,11)\n");
if(pixels_25_11!==16'h0051) $display("ERROR! at (25,11)\n");
if(pixels_26_11!==16'h070d) $display("ERROR! at (26,11)\n");
if(pixels_27_11!==16'h060e) $display("ERROR! at (27,11)\n");
if(pixels_28_11!==16'hfe18) $display("ERROR! at (28,11)\n");
if(pixels_29_11!==16'hfd3a) $display("ERROR! at (29,11)\n");
if(pixels_30_11!==16'h01e5) $display("ERROR! at (30,11)\n");
if(pixels_31_11!==16'hfff3) $display("ERROR! at (31,11)\n");
if(pixels_0_12!==16'hfeef) $display("ERROR! at (0,12)\n");
if(pixels_1_12!==16'h04e7) $display("ERROR! at (1,12)\n");
if(pixels_2_12!==16'h033a) $display("ERROR! at (2,12)\n");
if(pixels_3_12!==16'hf61e) $display("ERROR! at (3,12)\n");
if(pixels_4_12!==16'hff81) $display("ERROR! at (4,12)\n");
if(pixels_5_12!==16'h099a) $display("ERROR! at (5,12)\n");
if(pixels_6_12!==16'hfeaf) $display("ERROR! at (6,12)\n");
if(pixels_7_12!==16'hfb8d) $display("ERROR! at (7,12)\n");
if(pixels_8_12!==16'h0611) $display("ERROR! at (8,12)\n");
if(pixels_9_12!==16'hffc2) $display("ERROR! at (9,12)\n");
if(pixels_10_12!==16'hfbe6) $display("ERROR! at (10,12)\n");
if(pixels_11_12!==16'h0931) $display("ERROR! at (11,12)\n");
if(pixels_12_12!==16'hfc1e) $display("ERROR! at (12,12)\n");
if(pixels_13_12!==16'h014a) $display("ERROR! at (13,12)\n");
if(pixels_14_12!==16'hfe89) $display("ERROR! at (14,12)\n");
if(pixels_15_12!==16'hfb0c) $display("ERROR! at (15,12)\n");
if(pixels_16_12!==16'hfc61) $display("ERROR! at (16,12)\n");
if(pixels_17_12!==16'h0e47) $display("ERROR! at (17,12)\n");
if(pixels_18_12!==16'h07b7) $display("ERROR! at (18,12)\n");
if(pixels_19_12!==16'h05ee) $display("ERROR! at (19,12)\n");
if(pixels_20_12!==16'h026b) $display("ERROR! at (20,12)\n");
if(pixels_21_12!==16'hfe1c) $display("ERROR! at (21,12)\n");
if(pixels_22_12!==16'hf640) $display("ERROR! at (22,12)\n");
if(pixels_23_12!==16'h06c6) $display("ERROR! at (23,12)\n");
if(pixels_24_12!==16'h0500) $display("ERROR! at (24,12)\n");
if(pixels_25_12!==16'h00b2) $display("ERROR! at (25,12)\n");
if(pixels_26_12!==16'hffc9) $display("ERROR! at (26,12)\n");
if(pixels_27_12!==16'hfdc2) $display("ERROR! at (27,12)\n");
if(pixels_28_12!==16'h0527) $display("ERROR! at (28,12)\n");
if(pixels_29_12!==16'hfe56) $display("ERROR! at (29,12)\n");
if(pixels_30_12!==16'hfc3f) $display("ERROR! at (30,12)\n");
if(pixels_31_12!==16'hfc5e) $display("ERROR! at (31,12)\n");
if(pixels_0_13!==16'h022e) $display("ERROR! at (0,13)\n");
if(pixels_1_13!==16'h042f) $display("ERROR! at (1,13)\n");
if(pixels_2_13!==16'hfcdc) $display("ERROR! at (2,13)\n");
if(pixels_3_13!==16'hff60) $display("ERROR! at (3,13)\n");
if(pixels_4_13!==16'hff75) $display("ERROR! at (4,13)\n");
if(pixels_5_13!==16'hfa70) $display("ERROR! at (5,13)\n");
if(pixels_6_13!==16'hf8fa) $display("ERROR! at (6,13)\n");
if(pixels_7_13!==16'h01fb) $display("ERROR! at (7,13)\n");
if(pixels_8_13!==16'h0574) $display("ERROR! at (8,13)\n");
if(pixels_9_13!==16'hf9d4) $display("ERROR! at (9,13)\n");
if(pixels_10_13!==16'hf844) $display("ERROR! at (10,13)\n");
if(pixels_11_13!==16'hff51) $display("ERROR! at (11,13)\n");
if(pixels_12_13!==16'hf998) $display("ERROR! at (12,13)\n");
if(pixels_13_13!==16'h06b1) $display("ERROR! at (13,13)\n");
if(pixels_14_13!==16'h0717) $display("ERROR! at (14,13)\n");
if(pixels_15_13!==16'h02ff) $display("ERROR! at (15,13)\n");
if(pixels_16_13!==16'h05f0) $display("ERROR! at (16,13)\n");
if(pixels_17_13!==16'hffd2) $display("ERROR! at (17,13)\n");
if(pixels_18_13!==16'h03a1) $display("ERROR! at (18,13)\n");
if(pixels_19_13!==16'h0766) $display("ERROR! at (19,13)\n");
if(pixels_20_13!==16'hfc19) $display("ERROR! at (20,13)\n");
if(pixels_21_13!==16'hf89c) $display("ERROR! at (21,13)\n");
if(pixels_22_13!==16'hfa7f) $display("ERROR! at (22,13)\n");
if(pixels_23_13!==16'h000f) $display("ERROR! at (23,13)\n");
if(pixels_24_13!==16'h0021) $display("ERROR! at (24,13)\n");
if(pixels_25_13!==16'h0099) $display("ERROR! at (25,13)\n");
if(pixels_26_13!==16'hfd86) $display("ERROR! at (26,13)\n");
if(pixels_27_13!==16'hfe2a) $display("ERROR! at (27,13)\n");
if(pixels_28_13!==16'h001b) $display("ERROR! at (28,13)\n");
if(pixels_29_13!==16'h03fc) $display("ERROR! at (29,13)\n");
if(pixels_30_13!==16'h00b5) $display("ERROR! at (30,13)\n");
if(pixels_31_13!==16'hff99) $display("ERROR! at (31,13)\n");
if(pixels_0_14!==16'h0045) $display("ERROR! at (0,14)\n");
if(pixels_1_14!==16'hff31) $display("ERROR! at (1,14)\n");
if(pixels_2_14!==16'h0367) $display("ERROR! at (2,14)\n");
if(pixels_3_14!==16'hf5f2) $display("ERROR! at (3,14)\n");
if(pixels_4_14!==16'hfa6f) $display("ERROR! at (4,14)\n");
if(pixels_5_14!==16'h00b4) $display("ERROR! at (5,14)\n");
if(pixels_6_14!==16'hf4a2) $display("ERROR! at (6,14)\n");
if(pixels_7_14!==16'h00bd) $display("ERROR! at (7,14)\n");
if(pixels_8_14!==16'h02e8) $display("ERROR! at (8,14)\n");
if(pixels_9_14!==16'hfcf3) $display("ERROR! at (9,14)\n");
if(pixels_10_14!==16'h0545) $display("ERROR! at (10,14)\n");
if(pixels_11_14!==16'h039f) $display("ERROR! at (11,14)\n");
if(pixels_12_14!==16'hf8b8) $display("ERROR! at (12,14)\n");
if(pixels_13_14!==16'h0680) $display("ERROR! at (13,14)\n");
if(pixels_14_14!==16'hfed5) $display("ERROR! at (14,14)\n");
if(pixels_15_14!==16'hfb9b) $display("ERROR! at (15,14)\n");
if(pixels_16_14!==16'hfd70) $display("ERROR! at (16,14)\n");
if(pixels_17_14!==16'hffb2) $display("ERROR! at (17,14)\n");
if(pixels_18_14!==16'hf6f7) $display("ERROR! at (18,14)\n");
if(pixels_19_14!==16'hf113) $display("ERROR! at (19,14)\n");
if(pixels_20_14!==16'h0641) $display("ERROR! at (20,14)\n");
if(pixels_21_14!==16'hfd0f) $display("ERROR! at (21,14)\n");
if(pixels_22_14!==16'h003f) $display("ERROR! at (22,14)\n");
if(pixels_23_14!==16'hfa84) $display("ERROR! at (23,14)\n");
if(pixels_24_14!==16'h0081) $display("ERROR! at (24,14)\n");
if(pixels_25_14!==16'hfec7) $display("ERROR! at (25,14)\n");
if(pixels_26_14!==16'hffe9) $display("ERROR! at (26,14)\n");
if(pixels_27_14!==16'hf8e8) $display("ERROR! at (27,14)\n");
if(pixels_28_14!==16'h03fc) $display("ERROR! at (28,14)\n");
if(pixels_29_14!==16'h06b0) $display("ERROR! at (29,14)\n");
if(pixels_30_14!==16'h014f) $display("ERROR! at (30,14)\n");
if(pixels_31_14!==16'hfe44) $display("ERROR! at (31,14)\n");
if(pixels_0_15!==16'h0226) $display("ERROR! at (0,15)\n");
if(pixels_1_15!==16'h0414) $display("ERROR! at (1,15)\n");
if(pixels_2_15!==16'h0db1) $display("ERROR! at (2,15)\n");
if(pixels_3_15!==16'h0379) $display("ERROR! at (3,15)\n");
if(pixels_4_15!==16'hfdbf) $display("ERROR! at (4,15)\n");
if(pixels_5_15!==16'hfe1e) $display("ERROR! at (5,15)\n");
if(pixels_6_15!==16'h030a) $display("ERROR! at (6,15)\n");
if(pixels_7_15!==16'h1160) $display("ERROR! at (7,15)\n");
if(pixels_8_15!==16'hff8e) $display("ERROR! at (8,15)\n");
if(pixels_9_15!==16'h029f) $display("ERROR! at (9,15)\n");
if(pixels_10_15!==16'h022b) $display("ERROR! at (10,15)\n");
if(pixels_11_15!==16'hff96) $display("ERROR! at (11,15)\n");
if(pixels_12_15!==16'h0478) $display("ERROR! at (12,15)\n");
if(pixels_13_15!==16'h0377) $display("ERROR! at (13,15)\n");
if(pixels_14_15!==16'hf59a) $display("ERROR! at (14,15)\n");
if(pixels_15_15!==16'h05e8) $display("ERROR! at (15,15)\n");
if(pixels_16_15!==16'h04b3) $display("ERROR! at (16,15)\n");
if(pixels_17_15!==16'hf7e2) $display("ERROR! at (17,15)\n");
if(pixels_18_15!==16'hfaf0) $display("ERROR! at (18,15)\n");
if(pixels_19_15!==16'h02c2) $display("ERROR! at (19,15)\n");
if(pixels_20_15!==16'h0e3d) $display("ERROR! at (20,15)\n");
if(pixels_21_15!==16'hfe40) $display("ERROR! at (21,15)\n");
if(pixels_22_15!==16'h0a3d) $display("ERROR! at (22,15)\n");
if(pixels_23_15!==16'h000f) $display("ERROR! at (23,15)\n");
if(pixels_24_15!==16'hfda8) $display("ERROR! at (24,15)\n");
if(pixels_25_15!==16'h0646) $display("ERROR! at (25,15)\n");
if(pixels_26_15!==16'h02f4) $display("ERROR! at (26,15)\n");
if(pixels_27_15!==16'hfc4b) $display("ERROR! at (27,15)\n");
if(pixels_28_15!==16'h0036) $display("ERROR! at (28,15)\n");
if(pixels_29_15!==16'h0065) $display("ERROR! at (29,15)\n");
if(pixels_30_15!==16'hff10) $display("ERROR! at (30,15)\n");
if(pixels_31_15!==16'h0072) $display("ERROR! at (31,15)\n");
if(pixels_0_16!==16'h03fb) $display("ERROR! at (0,16)\n");
if(pixels_1_16!==16'h052d) $display("ERROR! at (1,16)\n");
if(pixels_2_16!==16'h051e) $display("ERROR! at (2,16)\n");
if(pixels_3_16!==16'hf81e) $display("ERROR! at (3,16)\n");
if(pixels_4_16!==16'hf911) $display("ERROR! at (4,16)\n");
if(pixels_5_16!==16'hfcf1) $display("ERROR! at (5,16)\n");
if(pixels_6_16!==16'hfd45) $display("ERROR! at (6,16)\n");
if(pixels_7_16!==16'h078f) $display("ERROR! at (7,16)\n");
if(pixels_8_16!==16'hf74c) $display("ERROR! at (8,16)\n");
if(pixels_9_16!==16'hf5dc) $display("ERROR! at (9,16)\n");
if(pixels_10_16!==16'hffb7) $display("ERROR! at (10,16)\n");
if(pixels_11_16!==16'h0bad) $display("ERROR! at (11,16)\n");
if(pixels_12_16!==16'h00ed) $display("ERROR! at (12,16)\n");
if(pixels_13_16!==16'hfbb9) $display("ERROR! at (13,16)\n");
if(pixels_14_16!==16'h019b) $display("ERROR! at (14,16)\n");
if(pixels_15_16!==16'h0fa3) $display("ERROR! at (15,16)\n");
if(pixels_16_16!==16'h0081) $display("ERROR! at (16,16)\n");
if(pixels_17_16!==16'hff6f) $display("ERROR! at (17,16)\n");
if(pixels_18_16!==16'h0b10) $display("ERROR! at (18,16)\n");
if(pixels_19_16!==16'h0812) $display("ERROR! at (19,16)\n");
if(pixels_20_16!==16'h0803) $display("ERROR! at (20,16)\n");
if(pixels_21_16!==16'hfdc6) $display("ERROR! at (21,16)\n");
if(pixels_22_16!==16'h0476) $display("ERROR! at (22,16)\n");
if(pixels_23_16!==16'hf98a) $display("ERROR! at (23,16)\n");
if(pixels_24_16!==16'hfba6) $display("ERROR! at (24,16)\n");
if(pixels_25_16!==16'h03a7) $display("ERROR! at (25,16)\n");
if(pixels_26_16!==16'hfc22) $display("ERROR! at (26,16)\n");
if(pixels_27_16!==16'hfc62) $display("ERROR! at (27,16)\n");
if(pixels_28_16!==16'hfcee) $display("ERROR! at (28,16)\n");
if(pixels_29_16!==16'hf9b8) $display("ERROR! at (29,16)\n");
if(pixels_30_16!==16'h01e2) $display("ERROR! at (30,16)\n");
if(pixels_31_16!==16'hfe02) $display("ERROR! at (31,16)\n");
if(pixels_0_17!==16'h00a2) $display("ERROR! at (0,17)\n");
if(pixels_1_17!==16'hff5b) $display("ERROR! at (1,17)\n");
if(pixels_2_17!==16'hfbdd) $display("ERROR! at (2,17)\n");
if(pixels_3_17!==16'h0352) $display("ERROR! at (3,17)\n");
if(pixels_4_17!==16'hfcf5) $display("ERROR! at (4,17)\n");
if(pixels_5_17!==16'h029f) $display("ERROR! at (5,17)\n");
if(pixels_6_17!==16'hf567) $display("ERROR! at (6,17)\n");
if(pixels_7_17!==16'hfecb) $display("ERROR! at (7,17)\n");
if(pixels_8_17!==16'hffd5) $display("ERROR! at (8,17)\n");
if(pixels_9_17!==16'h0581) $display("ERROR! at (9,17)\n");
if(pixels_10_17!==16'h04c4) $display("ERROR! at (10,17)\n");
if(pixels_11_17!==16'hfd3d) $display("ERROR! at (11,17)\n");
if(pixels_12_17!==16'hfe5d) $display("ERROR! at (12,17)\n");
if(pixels_13_17!==16'h007d) $display("ERROR! at (13,17)\n");
if(pixels_14_17!==16'h019e) $display("ERROR! at (14,17)\n");
if(pixels_15_17!==16'h0464) $display("ERROR! at (15,17)\n");
if(pixels_16_17!==16'hf9f1) $display("ERROR! at (16,17)\n");
if(pixels_17_17!==16'h0469) $display("ERROR! at (17,17)\n");
if(pixels_18_17!==16'hf8bc) $display("ERROR! at (18,17)\n");
if(pixels_19_17!==16'hf88f) $display("ERROR! at (19,17)\n");
if(pixels_20_17!==16'hf9f3) $display("ERROR! at (20,17)\n");
if(pixels_21_17!==16'hf9e0) $display("ERROR! at (21,17)\n");
if(pixels_22_17!==16'hf80c) $display("ERROR! at (22,17)\n");
if(pixels_23_17!==16'h02ff) $display("ERROR! at (23,17)\n");
if(pixels_24_17!==16'h073c) $display("ERROR! at (24,17)\n");
if(pixels_25_17!==16'hfe4f) $display("ERROR! at (25,17)\n");
if(pixels_26_17!==16'hfe1a) $display("ERROR! at (26,17)\n");
if(pixels_27_17!==16'h03ba) $display("ERROR! at (27,17)\n");
if(pixels_28_17!==16'h059a) $display("ERROR! at (28,17)\n");
if(pixels_29_17!==16'h04f3) $display("ERROR! at (29,17)\n");
if(pixels_30_17!==16'hffc8) $display("ERROR! at (30,17)\n");
if(pixels_31_17!==16'h033c) $display("ERROR! at (31,17)\n");
if(pixels_0_18!==16'h004a) $display("ERROR! at (0,18)\n");
if(pixels_1_18!==16'h0346) $display("ERROR! at (1,18)\n");
if(pixels_2_18!==16'h0121) $display("ERROR! at (2,18)\n");
if(pixels_3_18!==16'h0298) $display("ERROR! at (3,18)\n");
if(pixels_4_18!==16'h0ed1) $display("ERROR! at (4,18)\n");
if(pixels_5_18!==16'hfea8) $display("ERROR! at (5,18)\n");
if(pixels_6_18!==16'hfc15) $display("ERROR! at (6,18)\n");
if(pixels_7_18!==16'h03a8) $display("ERROR! at (7,18)\n");
if(pixels_8_18!==16'h0476) $display("ERROR! at (8,18)\n");
if(pixels_9_18!==16'hff21) $display("ERROR! at (9,18)\n");
if(pixels_10_18!==16'hff2f) $display("ERROR! at (10,18)\n");
if(pixels_11_18!==16'hfdd3) $display("ERROR! at (11,18)\n");
if(pixels_12_18!==16'hfa7d) $display("ERROR! at (12,18)\n");
if(pixels_13_18!==16'hff68) $display("ERROR! at (13,18)\n");
if(pixels_14_18!==16'hfd61) $display("ERROR! at (14,18)\n");
if(pixels_15_18!==16'hf810) $display("ERROR! at (15,18)\n");
if(pixels_16_18!==16'hf022) $display("ERROR! at (16,18)\n");
if(pixels_17_18!==16'h0179) $display("ERROR! at (17,18)\n");
if(pixels_18_18!==16'hfdee) $display("ERROR! at (18,18)\n");
if(pixels_19_18!==16'h03cb) $display("ERROR! at (19,18)\n");
if(pixels_20_18!==16'h0377) $display("ERROR! at (20,18)\n");
if(pixels_21_18!==16'hfe84) $display("ERROR! at (21,18)\n");
if(pixels_22_18!==16'h035b) $display("ERROR! at (22,18)\n");
if(pixels_23_18!==16'h0745) $display("ERROR! at (23,18)\n");
if(pixels_24_18!==16'hf5a6) $display("ERROR! at (24,18)\n");
if(pixels_25_18!==16'hfb74) $display("ERROR! at (25,18)\n");
if(pixels_26_18!==16'h02a5) $display("ERROR! at (26,18)\n");
if(pixels_27_18!==16'h01ed) $display("ERROR! at (27,18)\n");
if(pixels_28_18!==16'h0056) $display("ERROR! at (28,18)\n");
if(pixels_29_18!==16'hf8e2) $display("ERROR! at (29,18)\n");
if(pixels_30_18!==16'h0367) $display("ERROR! at (30,18)\n");
if(pixels_31_18!==16'h01cc) $display("ERROR! at (31,18)\n");
if(pixels_0_19!==16'hffb4) $display("ERROR! at (0,19)\n");
if(pixels_1_19!==16'hf918) $display("ERROR! at (1,19)\n");
if(pixels_2_19!==16'hf92f) $display("ERROR! at (2,19)\n");
if(pixels_3_19!==16'h080d) $display("ERROR! at (3,19)\n");
if(pixels_4_19!==16'h0119) $display("ERROR! at (4,19)\n");
if(pixels_5_19!==16'h007f) $display("ERROR! at (5,19)\n");
if(pixels_6_19!==16'hfd30) $display("ERROR! at (6,19)\n");
if(pixels_7_19!==16'hfb7b) $display("ERROR! at (7,19)\n");
if(pixels_8_19!==16'hfc49) $display("ERROR! at (8,19)\n");
if(pixels_9_19!==16'h0910) $display("ERROR! at (9,19)\n");
if(pixels_10_19!==16'h00be) $display("ERROR! at (10,19)\n");
if(pixels_11_19!==16'hfbc1) $display("ERROR! at (11,19)\n");
if(pixels_12_19!==16'h03c2) $display("ERROR! at (12,19)\n");
if(pixels_13_19!==16'h0cc1) $display("ERROR! at (13,19)\n");
if(pixels_14_19!==16'h0a00) $display("ERROR! at (14,19)\n");
if(pixels_15_19!==16'hf852) $display("ERROR! at (15,19)\n");
if(pixels_16_19!==16'hf4cc) $display("ERROR! at (16,19)\n");
if(pixels_17_19!==16'h0bca) $display("ERROR! at (17,19)\n");
if(pixels_18_19!==16'h03d8) $display("ERROR! at (18,19)\n");
if(pixels_19_19!==16'h01bf) $display("ERROR! at (19,19)\n");
if(pixels_20_19!==16'h0c27) $display("ERROR! at (20,19)\n");
if(pixels_21_19!==16'h0b6d) $display("ERROR! at (21,19)\n");
if(pixels_22_19!==16'h050e) $display("ERROR! at (22,19)\n");
if(pixels_23_19!==16'hfd6e) $display("ERROR! at (23,19)\n");
if(pixels_24_19!==16'hf747) $display("ERROR! at (24,19)\n");
if(pixels_25_19!==16'h0584) $display("ERROR! at (25,19)\n");
if(pixels_26_19!==16'h0626) $display("ERROR! at (26,19)\n");
if(pixels_27_19!==16'h0258) $display("ERROR! at (27,19)\n");
if(pixels_28_19!==16'hf9a7) $display("ERROR! at (28,19)\n");
if(pixels_29_19!==16'hfd8f) $display("ERROR! at (29,19)\n");
if(pixels_30_19!==16'hfa93) $display("ERROR! at (30,19)\n");
if(pixels_31_19!==16'hff99) $display("ERROR! at (31,19)\n");
if(pixels_0_20!==16'hfa7c) $display("ERROR! at (0,20)\n");
if(pixels_1_20!==16'hfe40) $display("ERROR! at (1,20)\n");
if(pixels_2_20!==16'h016f) $display("ERROR! at (2,20)\n");
if(pixels_3_20!==16'h00dd) $display("ERROR! at (3,20)\n");
if(pixels_4_20!==16'hff6e) $display("ERROR! at (4,20)\n");
if(pixels_5_20!==16'h02f5) $display("ERROR! at (5,20)\n");
if(pixels_6_20!==16'hfb05) $display("ERROR! at (6,20)\n");
if(pixels_7_20!==16'hf8a7) $display("ERROR! at (7,20)\n");
if(pixels_8_20!==16'h0828) $display("ERROR! at (8,20)\n");
if(pixels_9_20!==16'hfa25) $display("ERROR! at (9,20)\n");
if(pixels_10_20!==16'hff67) $display("ERROR! at (10,20)\n");
if(pixels_11_20!==16'h0142) $display("ERROR! at (11,20)\n");
if(pixels_12_20!==16'h0050) $display("ERROR! at (12,20)\n");
if(pixels_13_20!==16'h0d2a) $display("ERROR! at (13,20)\n");
if(pixels_14_20!==16'hfbae) $display("ERROR! at (14,20)\n");
if(pixels_15_20!==16'hf8ae) $display("ERROR! at (15,20)\n");
if(pixels_16_20!==16'h0462) $display("ERROR! at (16,20)\n");
if(pixels_17_20!==16'h029c) $display("ERROR! at (17,20)\n");
if(pixels_18_20!==16'hf8ef) $display("ERROR! at (18,20)\n");
if(pixels_19_20!==16'h015a) $display("ERROR! at (19,20)\n");
if(pixels_20_20!==16'h01a5) $display("ERROR! at (20,20)\n");
if(pixels_21_20!==16'hf8af) $display("ERROR! at (21,20)\n");
if(pixels_22_20!==16'hfb99) $display("ERROR! at (22,20)\n");
if(pixels_23_20!==16'hff54) $display("ERROR! at (23,20)\n");
if(pixels_24_20!==16'hf4fb) $display("ERROR! at (24,20)\n");
if(pixels_25_20!==16'h0549) $display("ERROR! at (25,20)\n");
if(pixels_26_20!==16'h0652) $display("ERROR! at (26,20)\n");
if(pixels_27_20!==16'h062a) $display("ERROR! at (27,20)\n");
if(pixels_28_20!==16'h06e3) $display("ERROR! at (28,20)\n");
if(pixels_29_20!==16'hfafa) $display("ERROR! at (29,20)\n");
if(pixels_30_20!==16'hff8b) $display("ERROR! at (30,20)\n");
if(pixels_31_20!==16'h03d4) $display("ERROR! at (31,20)\n");
if(pixels_0_21!==16'hfb96) $display("ERROR! at (0,21)\n");
if(pixels_1_21!==16'h05e9) $display("ERROR! at (1,21)\n");
if(pixels_2_21!==16'hfeef) $display("ERROR! at (2,21)\n");
if(pixels_3_21!==16'hff88) $display("ERROR! at (3,21)\n");
if(pixels_4_21!==16'h0426) $display("ERROR! at (4,21)\n");
if(pixels_5_21!==16'h069c) $display("ERROR! at (5,21)\n");
if(pixels_6_21!==16'hfc83) $display("ERROR! at (6,21)\n");
if(pixels_7_21!==16'h0352) $display("ERROR! at (7,21)\n");
if(pixels_8_21!==16'hf716) $display("ERROR! at (8,21)\n");
if(pixels_9_21!==16'h070a) $display("ERROR! at (9,21)\n");
if(pixels_10_21!==16'h0359) $display("ERROR! at (10,21)\n");
if(pixels_11_21!==16'hfee4) $display("ERROR! at (11,21)\n");
if(pixels_12_21!==16'hfa96) $display("ERROR! at (12,21)\n");
if(pixels_13_21!==16'hf5db) $display("ERROR! at (13,21)\n");
if(pixels_14_21!==16'hfaa0) $display("ERROR! at (14,21)\n");
if(pixels_15_21!==16'h0287) $display("ERROR! at (15,21)\n");
if(pixels_16_21!==16'hfe1b) $display("ERROR! at (16,21)\n");
if(pixels_17_21!==16'hf711) $display("ERROR! at (17,21)\n");
if(pixels_18_21!==16'hf899) $display("ERROR! at (18,21)\n");
if(pixels_19_21!==16'hf4b8) $display("ERROR! at (19,21)\n");
if(pixels_20_21!==16'hf96f) $display("ERROR! at (20,21)\n");
if(pixels_21_21!==16'h04b0) $display("ERROR! at (21,21)\n");
if(pixels_22_21!==16'h067d) $display("ERROR! at (22,21)\n");
if(pixels_23_21!==16'hfd2b) $display("ERROR! at (23,21)\n");
if(pixels_24_21!==16'hfa27) $display("ERROR! at (24,21)\n");
if(pixels_25_21!==16'hfedf) $display("ERROR! at (25,21)\n");
if(pixels_26_21!==16'h02dc) $display("ERROR! at (26,21)\n");
if(pixels_27_21!==16'hfffb) $display("ERROR! at (27,21)\n");
if(pixels_28_21!==16'hf89b) $display("ERROR! at (28,21)\n");
if(pixels_29_21!==16'hff78) $display("ERROR! at (29,21)\n");
if(pixels_30_21!==16'hfbe4) $display("ERROR! at (30,21)\n");
if(pixels_31_21!==16'hfcd6) $display("ERROR! at (31,21)\n");
if(pixels_0_22!==16'hff7d) $display("ERROR! at (0,22)\n");
if(pixels_1_22!==16'h099d) $display("ERROR! at (1,22)\n");
if(pixels_2_22!==16'hfbc2) $display("ERROR! at (2,22)\n");
if(pixels_3_22!==16'hf93e) $display("ERROR! at (3,22)\n");
if(pixels_4_22!==16'hf887) $display("ERROR! at (4,22)\n");
if(pixels_5_22!==16'hfcf6) $display("ERROR! at (5,22)\n");
if(pixels_6_22!==16'hffb5) $display("ERROR! at (6,22)\n");
if(pixels_7_22!==16'h012b) $display("ERROR! at (7,22)\n");
if(pixels_8_22!==16'hff80) $display("ERROR! at (8,22)\n");
if(pixels_9_22!==16'h02da) $display("ERROR! at (9,22)\n");
if(pixels_10_22!==16'h0387) $display("ERROR! at (10,22)\n");
if(pixels_11_22!==16'hfec0) $display("ERROR! at (11,22)\n");
if(pixels_12_22!==16'hfffa) $display("ERROR! at (12,22)\n");
if(pixels_13_22!==16'hfe63) $display("ERROR! at (13,22)\n");
if(pixels_14_22!==16'h03f3) $display("ERROR! at (14,22)\n");
if(pixels_15_22!==16'h0ae2) $display("ERROR! at (15,22)\n");
if(pixels_16_22!==16'h014d) $display("ERROR! at (16,22)\n");
if(pixels_17_22!==16'hff53) $display("ERROR! at (17,22)\n");
if(pixels_18_22!==16'hf8dd) $display("ERROR! at (18,22)\n");
if(pixels_19_22!==16'h0585) $display("ERROR! at (19,22)\n");
if(pixels_20_22!==16'h06a2) $display("ERROR! at (20,22)\n");
if(pixels_21_22!==16'h0763) $display("ERROR! at (21,22)\n");
if(pixels_22_22!==16'h033d) $display("ERROR! at (22,22)\n");
if(pixels_23_22!==16'h0d91) $display("ERROR! at (23,22)\n");
if(pixels_24_22!==16'hfd75) $display("ERROR! at (24,22)\n");
if(pixels_25_22!==16'h0086) $display("ERROR! at (25,22)\n");
if(pixels_26_22!==16'hf6d5) $display("ERROR! at (26,22)\n");
if(pixels_27_22!==16'h0504) $display("ERROR! at (27,22)\n");
if(pixels_28_22!==16'h0abb) $display("ERROR! at (28,22)\n");
if(pixels_29_22!==16'h04d9) $display("ERROR! at (29,22)\n");
if(pixels_30_22!==16'hfe43) $display("ERROR! at (30,22)\n");
if(pixels_31_22!==16'hfdcc) $display("ERROR! at (31,22)\n");
if(pixels_0_23!==16'h0043) $display("ERROR! at (0,23)\n");
if(pixels_1_23!==16'h01f1) $display("ERROR! at (1,23)\n");
if(pixels_2_23!==16'hf670) $display("ERROR! at (2,23)\n");
if(pixels_3_23!==16'hfd78) $display("ERROR! at (3,23)\n");
if(pixels_4_23!==16'h0219) $display("ERROR! at (4,23)\n");
if(pixels_5_23!==16'h00b2) $display("ERROR! at (5,23)\n");
if(pixels_6_23!==16'h01a9) $display("ERROR! at (6,23)\n");
if(pixels_7_23!==16'hfeb2) $display("ERROR! at (7,23)\n");
if(pixels_8_23!==16'hfb43) $display("ERROR! at (8,23)\n");
if(pixels_9_23!==16'h0019) $display("ERROR! at (9,23)\n");
if(pixels_10_23!==16'hfd1b) $display("ERROR! at (10,23)\n");
if(pixels_11_23!==16'h03d7) $display("ERROR! at (11,23)\n");
if(pixels_12_23!==16'hf768) $display("ERROR! at (12,23)\n");
if(pixels_13_23!==16'hff0b) $display("ERROR! at (13,23)\n");
if(pixels_14_23!==16'hffed) $display("ERROR! at (14,23)\n");
if(pixels_15_23!==16'hffc9) $display("ERROR! at (15,23)\n");
if(pixels_16_23!==16'hf9f7) $display("ERROR! at (16,23)\n");
if(pixels_17_23!==16'hf9b6) $display("ERROR! at (17,23)\n");
if(pixels_18_23!==16'h0416) $display("ERROR! at (18,23)\n");
if(pixels_19_23!==16'h07c7) $display("ERROR! at (19,23)\n");
if(pixels_20_23!==16'hf91c) $display("ERROR! at (20,23)\n");
if(pixels_21_23!==16'h02fe) $display("ERROR! at (21,23)\n");
if(pixels_22_23!==16'h042f) $display("ERROR! at (22,23)\n");
if(pixels_23_23!==16'h02ea) $display("ERROR! at (23,23)\n");
if(pixels_24_23!==16'hfb5e) $display("ERROR! at (24,23)\n");
if(pixels_25_23!==16'hfb93) $display("ERROR! at (25,23)\n");
if(pixels_26_23!==16'hfee4) $display("ERROR! at (26,23)\n");
if(pixels_27_23!==16'hf8b5) $display("ERROR! at (27,23)\n");
if(pixels_28_23!==16'h07ca) $display("ERROR! at (28,23)\n");
if(pixels_29_23!==16'h06d6) $display("ERROR! at (29,23)\n");
if(pixels_30_23!==16'h0223) $display("ERROR! at (30,23)\n");
if(pixels_31_23!==16'h0156) $display("ERROR! at (31,23)\n");
if(pixels_0_24!==16'hfee3) $display("ERROR! at (0,24)\n");
if(pixels_1_24!==16'hfbfd) $display("ERROR! at (1,24)\n");
if(pixels_2_24!==16'hff18) $display("ERROR! at (2,24)\n");
if(pixels_3_24!==16'h018e) $display("ERROR! at (3,24)\n");
if(pixels_4_24!==16'hfdcb) $display("ERROR! at (4,24)\n");
if(pixels_5_24!==16'hfabe) $display("ERROR! at (5,24)\n");
if(pixels_6_24!==16'h0042) $display("ERROR! at (6,24)\n");
if(pixels_7_24!==16'hff90) $display("ERROR! at (7,24)\n");
if(pixels_8_24!==16'h025f) $display("ERROR! at (8,24)\n");
if(pixels_9_24!==16'h0718) $display("ERROR! at (9,24)\n");
if(pixels_10_24!==16'hfb18) $display("ERROR! at (10,24)\n");
if(pixels_11_24!==16'h014b) $display("ERROR! at (11,24)\n");
if(pixels_12_24!==16'h031a) $display("ERROR! at (12,24)\n");
if(pixels_13_24!==16'hffe1) $display("ERROR! at (13,24)\n");
if(pixels_14_24!==16'hfd07) $display("ERROR! at (14,24)\n");
if(pixels_15_24!==16'h0083) $display("ERROR! at (15,24)\n");
if(pixels_16_24!==16'hfa42) $display("ERROR! at (16,24)\n");
if(pixels_17_24!==16'h013d) $display("ERROR! at (17,24)\n");
if(pixels_18_24!==16'h00c6) $display("ERROR! at (18,24)\n");
if(pixels_19_24!==16'hfc82) $display("ERROR! at (19,24)\n");
if(pixels_20_24!==16'hfea8) $display("ERROR! at (20,24)\n");
if(pixels_21_24!==16'hfd24) $display("ERROR! at (21,24)\n");
if(pixels_22_24!==16'hf469) $display("ERROR! at (22,24)\n");
if(pixels_23_24!==16'h0356) $display("ERROR! at (23,24)\n");
if(pixels_24_24!==16'hfd8a) $display("ERROR! at (24,24)\n");
if(pixels_25_24!==16'hfd69) $display("ERROR! at (25,24)\n");
if(pixels_26_24!==16'hfb3d) $display("ERROR! at (26,24)\n");
if(pixels_27_24!==16'h065e) $display("ERROR! at (27,24)\n");
if(pixels_28_24!==16'hff17) $display("ERROR! at (28,24)\n");
if(pixels_29_24!==16'hfc63) $display("ERROR! at (29,24)\n");
if(pixels_30_24!==16'hff02) $display("ERROR! at (30,24)\n");
if(pixels_31_24!==16'hfe24) $display("ERROR! at (31,24)\n");
if(pixels_0_25!==16'h01b9) $display("ERROR! at (0,25)\n");
if(pixels_1_25!==16'hff1c) $display("ERROR! at (1,25)\n");
if(pixels_2_25!==16'h036a) $display("ERROR! at (2,25)\n");
if(pixels_3_25!==16'h0c0b) $display("ERROR! at (3,25)\n");
if(pixels_4_25!==16'h0036) $display("ERROR! at (4,25)\n");
if(pixels_5_25!==16'h0084) $display("ERROR! at (5,25)\n");
if(pixels_6_25!==16'hfcdf) $display("ERROR! at (6,25)\n");
if(pixels_7_25!==16'hfae9) $display("ERROR! at (7,25)\n");
if(pixels_8_25!==16'hfd2f) $display("ERROR! at (8,25)\n");
if(pixels_9_25!==16'hfb50) $display("ERROR! at (9,25)\n");
if(pixels_10_25!==16'hf81a) $display("ERROR! at (10,25)\n");
if(pixels_11_25!==16'h0e0a) $display("ERROR! at (11,25)\n");
if(pixels_12_25!==16'h087c) $display("ERROR! at (12,25)\n");
if(pixels_13_25!==16'hffb3) $display("ERROR! at (13,25)\n");
if(pixels_14_25!==16'h05ab) $display("ERROR! at (14,25)\n");
if(pixels_15_25!==16'hfbb0) $display("ERROR! at (15,25)\n");
if(pixels_16_25!==16'hfe19) $display("ERROR! at (16,25)\n");
if(pixels_17_25!==16'hff83) $display("ERROR! at (17,25)\n");
if(pixels_18_25!==16'h02dd) $display("ERROR! at (18,25)\n");
if(pixels_19_25!==16'h0048) $display("ERROR! at (19,25)\n");
if(pixels_20_25!==16'h07a4) $display("ERROR! at (20,25)\n");
if(pixels_21_25!==16'h04d1) $display("ERROR! at (21,25)\n");
if(pixels_22_25!==16'hfbf8) $display("ERROR! at (22,25)\n");
if(pixels_23_25!==16'h055e) $display("ERROR! at (23,25)\n");
if(pixels_24_25!==16'hfef1) $display("ERROR! at (24,25)\n");
if(pixels_25_25!==16'h040a) $display("ERROR! at (25,25)\n");
if(pixels_26_25!==16'h0771) $display("ERROR! at (26,25)\n");
if(pixels_27_25!==16'hffcc) $display("ERROR! at (27,25)\n");
if(pixels_28_25!==16'hfa16) $display("ERROR! at (28,25)\n");
if(pixels_29_25!==16'hff64) $display("ERROR! at (29,25)\n");
if(pixels_30_25!==16'hfe79) $display("ERROR! at (30,25)\n");
if(pixels_31_25!==16'hfeb8) $display("ERROR! at (31,25)\n");
if(pixels_0_26!==16'h016d) $display("ERROR! at (0,26)\n");
if(pixels_1_26!==16'h0294) $display("ERROR! at (1,26)\n");
if(pixels_2_26!==16'h0099) $display("ERROR! at (2,26)\n");
if(pixels_3_26!==16'hfade) $display("ERROR! at (3,26)\n");
if(pixels_4_26!==16'hf7ad) $display("ERROR! at (4,26)\n");
if(pixels_5_26!==16'hff7c) $display("ERROR! at (5,26)\n");
if(pixels_6_26!==16'h00ff) $display("ERROR! at (6,26)\n");
if(pixels_7_26!==16'h0501) $display("ERROR! at (7,26)\n");
if(pixels_8_26!==16'h0350) $display("ERROR! at (8,26)\n");
if(pixels_9_26!==16'hfa78) $display("ERROR! at (9,26)\n");
if(pixels_10_26!==16'hfd6f) $display("ERROR! at (10,26)\n");
if(pixels_11_26!==16'h0632) $display("ERROR! at (11,26)\n");
if(pixels_12_26!==16'hfc0e) $display("ERROR! at (12,26)\n");
if(pixels_13_26!==16'h0737) $display("ERROR! at (13,26)\n");
if(pixels_14_26!==16'hf959) $display("ERROR! at (14,26)\n");
if(pixels_15_26!==16'hf7e9) $display("ERROR! at (15,26)\n");
if(pixels_16_26!==16'hfe3c) $display("ERROR! at (16,26)\n");
if(pixels_17_26!==16'h02d9) $display("ERROR! at (17,26)\n");
if(pixels_18_26!==16'hef5e) $display("ERROR! at (18,26)\n");
if(pixels_19_26!==16'hfd67) $display("ERROR! at (19,26)\n");
if(pixels_20_26!==16'hfa82) $display("ERROR! at (20,26)\n");
if(pixels_21_26!==16'hfc23) $display("ERROR! at (21,26)\n");
if(pixels_22_26!==16'h0043) $display("ERROR! at (22,26)\n");
if(pixels_23_26!==16'h05e7) $display("ERROR! at (23,26)\n");
if(pixels_24_26!==16'h04df) $display("ERROR! at (24,26)\n");
if(pixels_25_26!==16'h0511) $display("ERROR! at (25,26)\n");
if(pixels_26_26!==16'h0648) $display("ERROR! at (26,26)\n");
if(pixels_27_26!==16'hf827) $display("ERROR! at (27,26)\n");
if(pixels_28_26!==16'h0310) $display("ERROR! at (28,26)\n");
if(pixels_29_26!==16'h005c) $display("ERROR! at (29,26)\n");
if(pixels_30_26!==16'hff90) $display("ERROR! at (30,26)\n");
if(pixels_31_26!==16'h003a) $display("ERROR! at (31,26)\n");
if(pixels_0_27!==16'h0223) $display("ERROR! at (0,27)\n");
if(pixels_1_27!==16'hff3e) $display("ERROR! at (1,27)\n");
if(pixels_2_27!==16'h0253) $display("ERROR! at (2,27)\n");
if(pixels_3_27!==16'hfb3c) $display("ERROR! at (3,27)\n");
if(pixels_4_27!==16'hfced) $display("ERROR! at (4,27)\n");
if(pixels_5_27!==16'h0335) $display("ERROR! at (5,27)\n");
if(pixels_6_27!==16'hfdcb) $display("ERROR! at (6,27)\n");
if(pixels_7_27!==16'h02f8) $display("ERROR! at (7,27)\n");
if(pixels_8_27!==16'h017c) $display("ERROR! at (8,27)\n");
if(pixels_9_27!==16'hfeb2) $display("ERROR! at (9,27)\n");
if(pixels_10_27!==16'h02c5) $display("ERROR! at (10,27)\n");
if(pixels_11_27!==16'h08f2) $display("ERROR! at (11,27)\n");
if(pixels_12_27!==16'hfcc4) $display("ERROR! at (12,27)\n");
if(pixels_13_27!==16'hfd46) $display("ERROR! at (13,27)\n");
if(pixels_14_27!==16'hfd50) $display("ERROR! at (14,27)\n");
if(pixels_15_27!==16'h0a52) $display("ERROR! at (15,27)\n");
if(pixels_16_27!==16'h0477) $display("ERROR! at (16,27)\n");
if(pixels_17_27!==16'hfdd2) $display("ERROR! at (17,27)\n");
if(pixels_18_27!==16'h095c) $display("ERROR! at (18,27)\n");
if(pixels_19_27!==16'h0089) $display("ERROR! at (19,27)\n");
if(pixels_20_27!==16'hff61) $display("ERROR! at (20,27)\n");
if(pixels_21_27!==16'h002b) $display("ERROR! at (21,27)\n");
if(pixels_22_27!==16'h0663) $display("ERROR! at (22,27)\n");
if(pixels_23_27!==16'h00cd) $display("ERROR! at (23,27)\n");
if(pixels_24_27!==16'h067e) $display("ERROR! at (24,27)\n");
if(pixels_25_27!==16'h0328) $display("ERROR! at (25,27)\n");
if(pixels_26_27!==16'hf6d1) $display("ERROR! at (26,27)\n");
if(pixels_27_27!==16'hf8c5) $display("ERROR! at (27,27)\n");
if(pixels_28_27!==16'h0654) $display("ERROR! at (28,27)\n");
if(pixels_29_27!==16'h02ca) $display("ERROR! at (29,27)\n");
if(pixels_30_27!==16'h015c) $display("ERROR! at (30,27)\n");
if(pixels_31_27!==16'hff7d) $display("ERROR! at (31,27)\n");
if(pixels_0_28!==16'h012c) $display("ERROR! at (0,28)\n");
if(pixels_1_28!==16'hfc9f) $display("ERROR! at (1,28)\n");
if(pixels_2_28!==16'h051e) $display("ERROR! at (2,28)\n");
if(pixels_3_28!==16'h030e) $display("ERROR! at (3,28)\n");
if(pixels_4_28!==16'h025e) $display("ERROR! at (4,28)\n");
if(pixels_5_28!==16'h0429) $display("ERROR! at (5,28)\n");
if(pixels_6_28!==16'hfacb) $display("ERROR! at (6,28)\n");
if(pixels_7_28!==16'hfeac) $display("ERROR! at (7,28)\n");
if(pixels_8_28!==16'hfcec) $display("ERROR! at (8,28)\n");
if(pixels_9_28!==16'hfdd8) $display("ERROR! at (9,28)\n");
if(pixels_10_28!==16'h0037) $display("ERROR! at (10,28)\n");
if(pixels_11_28!==16'h0593) $display("ERROR! at (11,28)\n");
if(pixels_12_28!==16'hf9b8) $display("ERROR! at (12,28)\n");
if(pixels_13_28!==16'h0152) $display("ERROR! at (13,28)\n");
if(pixels_14_28!==16'h08bd) $display("ERROR! at (14,28)\n");
if(pixels_15_28!==16'hff93) $display("ERROR! at (15,28)\n");
if(pixels_16_28!==16'hfb44) $display("ERROR! at (16,28)\n");
if(pixels_17_28!==16'h05bc) $display("ERROR! at (17,28)\n");
if(pixels_18_28!==16'hfbf7) $display("ERROR! at (18,28)\n");
if(pixels_19_28!==16'hf812) $display("ERROR! at (19,28)\n");
if(pixels_20_28!==16'hfdb9) $display("ERROR! at (20,28)\n");
if(pixels_21_28!==16'h0008) $display("ERROR! at (21,28)\n");
if(pixels_22_28!==16'h026f) $display("ERROR! at (22,28)\n");
if(pixels_23_28!==16'h02a3) $display("ERROR! at (23,28)\n");
if(pixels_24_28!==16'h0912) $display("ERROR! at (24,28)\n");
if(pixels_25_28!==16'hf89a) $display("ERROR! at (25,28)\n");
if(pixels_26_28!==16'hfe66) $display("ERROR! at (26,28)\n");
if(pixels_27_28!==16'h00d5) $display("ERROR! at (27,28)\n");
if(pixels_28_28!==16'hfd7a) $display("ERROR! at (28,28)\n");
if(pixels_29_28!==16'h0078) $display("ERROR! at (29,28)\n");
if(pixels_30_28!==16'hfe6e) $display("ERROR! at (30,28)\n");
if(pixels_31_28!==16'hff28) $display("ERROR! at (31,28)\n");
if(pixels_0_29!==16'hffd9) $display("ERROR! at (0,29)\n");
if(pixels_1_29!==16'hfe9f) $display("ERROR! at (1,29)\n");
if(pixels_2_29!==16'h0150) $display("ERROR! at (2,29)\n");
if(pixels_3_29!==16'hff5f) $display("ERROR! at (3,29)\n");
if(pixels_4_29!==16'h03f0) $display("ERROR! at (4,29)\n");
if(pixels_5_29!==16'hfe25) $display("ERROR! at (5,29)\n");
if(pixels_6_29!==16'hfc90) $display("ERROR! at (6,29)\n");
if(pixels_7_29!==16'hfe1a) $display("ERROR! at (7,29)\n");
if(pixels_8_29!==16'hfdf3) $display("ERROR! at (8,29)\n");
if(pixels_9_29!==16'hfe94) $display("ERROR! at (9,29)\n");
if(pixels_10_29!==16'h00ed) $display("ERROR! at (10,29)\n");
if(pixels_11_29!==16'hffdd) $display("ERROR! at (11,29)\n");
if(pixels_12_29!==16'hfe2b) $display("ERROR! at (12,29)\n");
if(pixels_13_29!==16'h04c2) $display("ERROR! at (13,29)\n");
if(pixels_14_29!==16'hfff2) $display("ERROR! at (14,29)\n");
if(pixels_15_29!==16'hfefe) $display("ERROR! at (15,29)\n");
if(pixels_16_29!==16'hffa6) $display("ERROR! at (16,29)\n");
if(pixels_17_29!==16'hfb4d) $display("ERROR! at (17,29)\n");
if(pixels_18_29!==16'hfdba) $display("ERROR! at (18,29)\n");
if(pixels_19_29!==16'hfee5) $display("ERROR! at (19,29)\n");
if(pixels_20_29!==16'hfd75) $display("ERROR! at (20,29)\n");
if(pixels_21_29!==16'hfa45) $display("ERROR! at (21,29)\n");
if(pixels_22_29!==16'hfb4c) $display("ERROR! at (22,29)\n");
if(pixels_23_29!==16'hf9e2) $display("ERROR! at (23,29)\n");
if(pixels_24_29!==16'hffb6) $display("ERROR! at (24,29)\n");
if(pixels_25_29!==16'h00d0) $display("ERROR! at (25,29)\n");
if(pixels_26_29!==16'h0631) $display("ERROR! at (26,29)\n");
if(pixels_27_29!==16'hfff1) $display("ERROR! at (27,29)\n");
if(pixels_28_29!==16'h02e0) $display("ERROR! at (28,29)\n");
if(pixels_29_29!==16'hfe5e) $display("ERROR! at (29,29)\n");
if(pixels_30_29!==16'hfe07) $display("ERROR! at (30,29)\n");
if(pixels_31_29!==16'hfff3) $display("ERROR! at (31,29)\n");
if(pixels_0_30!==16'hffc3) $display("ERROR! at (0,30)\n");
if(pixels_1_30!==16'h0067) $display("ERROR! at (1,30)\n");
if(pixels_2_30!==16'hffba) $display("ERROR! at (2,30)\n");
if(pixels_3_30!==16'hfff8) $display("ERROR! at (3,30)\n");
if(pixels_4_30!==16'h009b) $display("ERROR! at (4,30)\n");
if(pixels_5_30!==16'h00ea) $display("ERROR! at (5,30)\n");
if(pixels_6_30!==16'h00ce) $display("ERROR! at (6,30)\n");
if(pixels_7_30!==16'h0381) $display("ERROR! at (7,30)\n");
if(pixels_8_30!==16'h02b8) $display("ERROR! at (8,30)\n");
if(pixels_9_30!==16'h0020) $display("ERROR! at (9,30)\n");
if(pixels_10_30!==16'h00d0) $display("ERROR! at (10,30)\n");
if(pixels_11_30!==16'hfd8a) $display("ERROR! at (11,30)\n");
if(pixels_12_30!==16'hff92) $display("ERROR! at (12,30)\n");
if(pixels_13_30!==16'h0221) $display("ERROR! at (13,30)\n");
if(pixels_14_30!==16'h02f9) $display("ERROR! at (14,30)\n");
if(pixels_15_30!==16'hfe16) $display("ERROR! at (15,30)\n");
if(pixels_16_30!==16'h020b) $display("ERROR! at (16,30)\n");
if(pixels_17_30!==16'h0441) $display("ERROR! at (17,30)\n");
if(pixels_18_30!==16'h044b) $display("ERROR! at (18,30)\n");
if(pixels_19_30!==16'h01a3) $display("ERROR! at (19,30)\n");
if(pixels_20_30!==16'h055e) $display("ERROR! at (20,30)\n");
if(pixels_21_30!==16'h02d0) $display("ERROR! at (21,30)\n");
if(pixels_22_30!==16'hffdf) $display("ERROR! at (22,30)\n");
if(pixels_23_30!==16'h0048) $display("ERROR! at (23,30)\n");
if(pixels_24_30!==16'hffec) $display("ERROR! at (24,30)\n");
if(pixels_25_30!==16'h012e) $display("ERROR! at (25,30)\n");
if(pixels_26_30!==16'h0273) $display("ERROR! at (26,30)\n");
if(pixels_27_30!==16'h0300) $display("ERROR! at (27,30)\n");
if(pixels_28_30!==16'hfd6e) $display("ERROR! at (28,30)\n");
if(pixels_29_30!==16'hff49) $display("ERROR! at (29,30)\n");
if(pixels_30_30!==16'h00bb) $display("ERROR! at (30,30)\n");
if(pixels_31_30!==16'h00a6) $display("ERROR! at (31,30)\n");
if(pixels_0_31!==16'hffb8) $display("ERROR! at (0,31)\n");
if(pixels_1_31!==16'h0090) $display("ERROR! at (1,31)\n");
if(pixels_2_31!==16'hffd2) $display("ERROR! at (2,31)\n");
if(pixels_3_31!==16'hff24) $display("ERROR! at (3,31)\n");
if(pixels_4_31!==16'hff98) $display("ERROR! at (4,31)\n");
if(pixels_5_31!==16'h00de) $display("ERROR! at (5,31)\n");
if(pixels_6_31!==16'hff4a) $display("ERROR! at (6,31)\n");
if(pixels_7_31!==16'h005c) $display("ERROR! at (7,31)\n");
if(pixels_8_31!==16'hff40) $display("ERROR! at (8,31)\n");
if(pixels_9_31!==16'hfecc) $display("ERROR! at (9,31)\n");
if(pixels_10_31!==16'hfffa) $display("ERROR! at (10,31)\n");
if(pixels_11_31!==16'hfee0) $display("ERROR! at (11,31)\n");
if(pixels_12_31!==16'h002e) $display("ERROR! at (12,31)\n");
if(pixels_13_31!==16'h013a) $display("ERROR! at (13,31)\n");
if(pixels_14_31!==16'hff86) $display("ERROR! at (14,31)\n");
if(pixels_15_31!==16'hfda6) $display("ERROR! at (15,31)\n");
if(pixels_16_31!==16'h0168) $display("ERROR! at (16,31)\n");
if(pixels_17_31!==16'hff7a) $display("ERROR! at (17,31)\n");
if(pixels_18_31!==16'hfd6c) $display("ERROR! at (18,31)\n");
if(pixels_19_31!==16'hfffa) $display("ERROR! at (19,31)\n");
if(pixels_20_31!==16'h006e) $display("ERROR! at (20,31)\n");
if(pixels_21_31!==16'hfe8e) $display("ERROR! at (21,31)\n");
if(pixels_22_31!==16'hfe6a) $display("ERROR! at (22,31)\n");
if(pixels_23_31!==16'hffe4) $display("ERROR! at (23,31)\n");
if(pixels_24_31!==16'hfe8a) $display("ERROR! at (24,31)\n");
if(pixels_25_31!==16'h00f4) $display("ERROR! at (25,31)\n");
if(pixels_26_31!==16'h015e) $display("ERROR! at (26,31)\n");
if(pixels_27_31!==16'hff6e) $display("ERROR! at (27,31)\n");
if(pixels_28_31!==16'hfde4) $display("ERROR! at (28,31)\n");
if(pixels_29_31!==16'h0136) $display("ERROR! at (29,31)\n");
if(pixels_30_31!==16'hff5e) $display("ERROR! at (30,31)\n");
if(pixels_31_31!==16'hffb8) $display("ERROR! at (31,31)\n");





    $finish;

end

always@(posedge clk)begin
    if(out_valid)begin
        
        result[ (($signed(col_answer_1_1)+4)+($signed(row_answer_1_1)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_1_1)+4)+($signed(row_answer_1_1)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_1_1);
        result[ (($signed(col_answer_1_2)+4)+($signed(row_answer_1_2)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_1_2)+4)+($signed(row_answer_1_2)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_1_2);
        result[ (($signed(col_answer_1_3)+4)+($signed(row_answer_1_3)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_1_3)+4)+($signed(row_answer_1_3)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_1_3);
        result[ (($signed(col_answer_1_4)+4)+($signed(row_answer_1_4)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_1_4)+4)+($signed(row_answer_1_4)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_1_4);

        result[ (($signed(col_answer_2_1)+4)+($signed(row_answer_2_1)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_2_1)+4)+($signed(row_answer_2_1)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_2_1);
        result[ (($signed(col_answer_2_2)+4)+($signed(row_answer_2_2)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_2_2)+4)+($signed(row_answer_2_2)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_2_2);
        result[ (($signed(col_answer_2_3)+4)+($signed(row_answer_2_3)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_2_3)+4)+($signed(row_answer_2_3)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_2_3);
        result[ (($signed(col_answer_2_4)+4)+($signed(row_answer_2_4)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_2_4)+4)+($signed(row_answer_2_4)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_2_4);

        result[ (($signed(col_answer_3_1)+4)+($signed(row_answer_3_1)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_3_1)+4)+($signed(row_answer_3_1)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_3_1);
        result[ (($signed(col_answer_3_2)+4)+($signed(row_answer_3_2)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_3_2)+4)+($signed(row_answer_3_2)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_3_2);
        result[ (($signed(col_answer_3_3)+4)+($signed(row_answer_3_3)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_3_3)+4)+($signed(row_answer_3_3)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_3_3);
        result[ (($signed(col_answer_3_4)+4)+($signed(row_answer_3_4)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_3_4)+4)+($signed(row_answer_3_4)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_3_4);

        result[ (($signed(col_answer_4_1)+4)+($signed(row_answer_4_1)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_4_1)+4)+($signed(row_answer_4_1)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_4_1);
        result[ (($signed(col_answer_4_2)+4)+($signed(row_answer_4_2)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_4_2)+4)+($signed(row_answer_4_2)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_4_2);
        result[ (($signed(col_answer_4_3)+4)+($signed(row_answer_4_3)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_4_3)+4)+($signed(row_answer_4_3)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_4_3);
        result[ (($signed(col_answer_4_4)+4)+($signed(row_answer_4_4)+4)*32+1)*word_length*2-1 -:word_length*2] = $signed(result[ (($signed(col_answer_4_4)+4)+($signed(row_answer_4_4)+4)*32+1)*word_length*2-1 -:word_length*2]) + $signed(answer_4_4);

    end
    //result[11*(data_out_rows[col_length-1:0]+4)+(data_out_cols[col_length-1:0]+4)+1 -:word_length] <= data_out[word_length-1:0] + result[11*(data_out_rows[col_length-1:0]+4)+(data_out_cols[col_length-1:0]+4)+1 -:word_length];
end


always #5 clk = ~clk;




PE #(
    .col_length(col_length), 
    .word_length(word_length), 
    .double_word_length(double_word_length), 
    .kernel_size(kernel_size), 
    .image_size(image_size)
    ) pe_TOP( 
    .clk(clk), 
    .rst(rst), 
    .in_valid(in_valid),
    .feature_valid_num(feature_valid_num),
    .feature_value(pe_input_feature_value),
    .feature_cols(pe_input_feature_cols),
    .feature_rows(pe_input_feature_rows),
    .weight_valid_num(weight_valid_num),
    .weight_value(pe_input_weight_value),
    .weight_cols(pe_input_weight_cols),
    .weight_rows(pe_input_weight_rows),
    .data_out(data_out),
    .data_out_cols(data_out_cols),
    .data_out_rows(data_out_rows),
    .out_valid(out_valid)
);







endmodule